--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--#CCDOF0HMCR#0CR8VHHM0MHF3WRRCHRIDCDRP0CMkDND$8RN8DRLF_O	sRFl0
FF-N-RsDOEHR#0=CR#D0CO_lsF

---f-R]8CNCRs:/$/#MHbDO$H0/blNolI/NCbbsG#/HMDHGH/DLC/oMHCsOC/oMC_oMHCsOF/slE3P8Ry4f-
-
H
DLssN$CRHC
C;
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RsIF	C3oMObN	CNo3DND;D

HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00)$RmLv_NR#CHS#
oCCMsRHO5S
SS8IH0:ERR0HMCsoCRR:=cS;
S8SN8HsI8R0E:MRH0CCos=R:R
(;SDSSF8IN8:sRR0HMCsoCRR:=jS;
SHSEo8EN8:sRR0HMCsoCRR:=(
U;S0SSNCLDRs:RFNl0L;DC
SSS80VDRs:RFFlIsS8
2S;
b0FsRS5
S7Sq7:)RRRHM#_08DHFoOC_POs0FR85N8HsI8R0E-RR48MFI0jFR2S;
SmS7z:aRR0FkR8#0_oDFHPO_CFO0sIR5HE80R4-RRI8FMR0FjS2
S
2;S0N0skHL0QCRhRQa:0R#soHM;N
S0H0sLCk0Rs\3N\M	RH:RMo0CC
s;RRRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MC8RM00H$mR)vN_L#
C;
ONsECH0Os0kCCR#D0CO_v)mRRFV)_mvLCN#R
H#SL#k0C$bRlsFFRk0H##R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2-;
-FSOlMbFCRM0vwzXn-
-SFSbs50R
S--SmSSRRR:FRk0#_08DHFoO-;
-SSSSRQj:MRHR8#0_oDFH
O;-S-SS4SQRH:RM0R#8F_Do;HO
S--S1SSRRR:H#MR0D8_FOoH
S--S;S2
S--CRM8ObFlFMMC0
;S
FSOMN#0ME0RC:GRRs#0H5MojFR0R246RR:=".j4dnc6(qUgA B7w
";
kSVMHO0FsMRFNl0LsDCC5N80DNLCRR:s0FlNCLD;,RIRRL,DRCM:MRH0CCoss2RCs0kM0R#soHMRR=>"lsF0DNLCNsC8
";
kSVMHO0FVMRkPMONLD5FF00lMDHC,_VRIDFNs88_RV,EEHoNs88_RV,L,H0RHML0:#RR0HMCsoC2CRs0MksRs#0HRMoHS#
SMOF#M0N0FR0bRR:HCM0oRCs:L=RFF00lMDHCR_V+LRMHR0#-;R4
PSSNNsHLRDCH[,R,,RPRFLb#RR:HCM0o;Cs
OSSF0M#NRM00OFbERNs:MRH0CCos=R:RHML0/#RR-cRR
4;SNSPsLHNDLCRk:VRRs#0H5Mo0OFbERNs8MFI0jFR2S;
LHCoMS
SHLV5FF00lMDHCR_V<FRDI8N8sR_VF0sRF>bRRoEHE8N8s2_VRC0EMS
SS:[R=;Rj
SSSP=R:R
j;SLSSbRF#:j=R;S
SSsVFRHHRMFRL0l0FDCHM_0VRFFR0bDRRF
FbSSSSHHVRRD<RF8IN8Vs_RRFsHRR>EEHoNs88_0VRE
CMSSSSSRHV80VD50LH2RR='R4'0MEC
SSSSPSSRR:=PRR+.[**;S
SSCSSMH8RVS;
SCSSD
#CSSSSSRHV0DNLC25H50LH2RR='R4'0MEC
SSSSPSSRR:=PRR+.[**;S
SSCSSMH8RVS;
SCSSMH8RVS;
S[SSRR:=[RR+4R;RR-R-RlMkLRCsFLVRHR0#ODFDCCO08SR
SHSSVR5[=2RcRC0EM-R-RCCPsc$RRRIC8bklR0HMFRRNOsENNCO0sS
SS[SSRR:=jS;
SSSSL5kVL#bF2=R:RGEC5;P2
SSSSbSLF:#R=bRLF+#RR
4;SSSSS:PR=;Rj
SSSS8CMR;HV
SSSCRM8DbFF;S
SS0sCkRsML;kV
CSSD
#CSsSSCs0kMFRslL0NDCCsN085NCLD,FRL0l0FDCHM_RV,L,H0RHML0;#2
CSSMH8RVS;
CRM8VOkM0MHFRMVkODPN;S

O#FM00NMR0LF0pFlHRMC:MRH0CCos=R:RF5DI8N8sn/42n*4;O
SF0M#NRM0L0F0F.ldpCHMRH:RMo0CC:sR=DR5F8IN8ds/.d2*.S;
O#FM00NMRoEHEMpHCRR:HCM0oRCs:5=REEHoNs88/24n*;4n
FSOMN#0ME0RHdoE.MpHCRR:HCM0oRCs:5=REEHoNs88/2d.*;d.
FSOMN#0ME0RHAoEFCs8sRR:HCM0oRCs:E=RHpoEHRMC+6R4RS;
O#FM00NMRH0s#00NCR_H:MRH0CCos=R:RH5EoFEAss8C+L4-FF00lMpHC42/n
R;Sb0$CNR0L#RHRsNsN5$R5oEHEpd.HRMC-FRL0l0FdH.pM/C2d4.+RI8FMR0FjF2RVFRsl0FkRS;
#MHoN1DRm,zaRzpmaRR:0;NL
HS#oDMNRz7mak_NG7,Rm_zaN.kGR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2L;
CMoH
RRRRFRVsH_bbRC:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0SC
S0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#;R4
RRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoRD:RNDLCRRH#4S;
RoLCHSM
SCRsoR#:bCHbL
kVSRSSb0FsRblN5R
SRSRSSRSRQ>R=Rz7mak_NG25H,R
SRSRSSRSRm>R=Rz7ma25H
SSSS2SR;R
SCRM8oCCMsCN0RsVF_bbHC
;
S_HV4:n#RRHV5oEHEpd.HRMC>FRL0l0FdH.pMRC2oCCMsCN0
LSSCMoH
HSSVn_4LH:RVLR5FF00lMpHCRR=L0F0F.ldpCHM2CRoMNCs0SC
S:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSSSSNs00H0LkChRQQFaRVmR)vR 6:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL0d,R.
2;SLSSCMoH
SSSSv)m :6RRv)md4.X
SSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSqSS4>R=R7q7)254,S
SSSSSSqSS.>R=R7q7)25.,S
SSSSSSqSSd>R=R7q7)25d,S
SSSSSSqSSc>R=R7q7)25c,S
SSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SS8CMRMoCC0sNC;RL
CSSMo8RCsMCNR0CH4V_n
L;SVSH_L4n:VRHRF5L0l0FpCHMRL>RFF00lpd.H2MCRMoCC0sNCS
SSRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SNSS0H0sLCk0RQQhaVRFRv)m :cRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SCSLo
HMSSSS) mvcRR:)4mvn
X4SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSS4SqRR=>q)775,42
SSSSSSSS.SqRR=>q)775,.2
SSSSSSSSdSqRR=>q)775,d2
SSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSCRM8oCCMsCN0R
L;SMSC8CRoMNCs0HCRVn_4LS;
CRM8oCCMsCN0R_HV4;n#
H
SV._d#H:RVER5HdoE.MpHCRR=L0F0F.ldpCHM2CRoMNCs0SC
S_HV4:nORRHV50LF0pFlHRMC=FRL0l0FdH.pMRC2oCCMsCN0
SSSLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SSVSH_R4:H5VRNs88I0H8ERR=4o2RCsMCN
0CSSSSS0N0skHL0QCRhRQaF)VRm4v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSoLCHSM
SSSS) mv4RR:)4mvn
X4SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSq=4R>jR''S,
SSSSSSSSSRq.='>Rj
',SSSSSSSSSdSqRR=>',j'
SSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SSMSC8CRoMNCs0HCRV;_4
SSSS_HV.H:RVNR58I8sHE80R.=R2CRoMNCs0SC
SSSSNs00H0LkChRQQFaRVmR)vR .:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSLHCoMS
SS)SSm.v R):Rmnv4XS4
SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSq=.R>jR''S,
SSSSSSSSSRqd='>Rj
',SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSS8CMRMoCC0sNCVRH_
.;SSSSHdV_:VRHR85N8HsI8R0E=2RdRMoCC0sNCS
SSNSS0H0sLCk0RQQhaVRFRv)m :dRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SLSSCMoH
SSSSmS)vR d:mR)vX4n4S
SSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSq=dR>jR''S,
SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSS2SS;S
SSMSC8CRoMNCs0HCRV;_d
SSSS_HVcH:RV5R5EEHoNs88-0LF0pFlHRMC<nR42MRN8NR58I8sHE80RR>=cR22oCCMsCN0
SSSS0SN0LsHkR0CQahQRRFV) mvcRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSCSLo
HMSSSSSv)m :cRRv)m44nX
SSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSqSSd>R=R7q7)25d,S
SSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SCSSMo8RCsMCNR0CHcV_;S
SSVSH_R6:H5VR58N8s8IH0>ER=2R6R8NMRH5Eo8EN8-sRR0LF0pFlHRMC>4=RnR22oCCMsCN0
SSSS0SN0LsHkR0CQahQRRFV) mv6RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R2d.;S
SSCSLo
HMSSSSSv)m :6RRv)md4.X
SSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSSRq4=q>R757)4
2,SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSqSSd>R=R7q7)25d,S
SSSSSSSSSq=cR>7Rq7c)52S,
SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SSSSCRM8oCCMsCN0R_HV6S;
SMSC8CRoMNCs0LCR;S
SCRM8oCCMsCN0R_HV4;nO
HSSVn_48H:RVLR5FF00lMpHCRR>L0F0F.ldpCHM2CRoMNCs0SC
SVSH_sN8I0H8EH:RVNR58I8sHE80Rc>R2CRoMNCs0SC
SLSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSSVSH_Rc:H5VR5oEHE8N8sF-L0l0FDCHMR4<RnN2RM58RNs88I0H8E=R>R2c2RMoCC0sNCS
SSSSSNs00H0LkChRQQFaRVmR)vR c:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSSoLCHSM
SSSSSv)m :cRRv)m44nX
SSSSSSSSsbF0NRlbRR5q=jR>7Rq7j)52S,
SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSdSqRR=>q)775,d2
SSSSSSSSSSSm>R=Rz1ma25j50LH2S
SSSSSSSSSS
2;SSSSS8CMRMoCC0sNCVRH_
c;SSSSCRM8oCCMsCN0R
L;SCSSMo8RCsMCNR0CHNV_8HsI8;0E
SSSHNV_8I8sHE80:VRHR85N8HsI8R0E<c=R2CRoMNCs0SC
SLSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSSVSH_R4:H5VRNs88I0H8ERR=4o2RCsMCN
0CSSSSS0SN0LsHkR0CQahQRRFV) mv4RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSLSSCMoH
SSSS)SSm4v R):Rmnv4XS4
SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSSRq4='>Rj
',SSSSSSSSSqSS.>R=R''j,S
SSSSSSSSSSRqd='>Rj
',SSSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSSSSS2S;
SSSSCRM8oCCMsCN0R_HV4S;
SSSSH.V_:VRHR85N8HsI8R0E=2R.RMoCC0sNCS
SSSSSNs00H0LkChRQQFaRVmR)vR .:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSSoLCHSM
SSSSSv)m :.RRv)m44nX
SSSSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSSRq.='>Rj
',SSSSSSSSSqSSd>R=R''j,S
SSSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS;S2
SSSSMSC8CRoMNCs0HCRV;_.
SSSSVSH_Rd:H5VRNs88I0H8ERR=do2RCsMCN
0CSSSSS0SN0LsHkR0CQahQRRFV) mvdRR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSLSSCMoH
SSSS)SSmdv R):Rmnv4XS4
SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSSRq4=q>R757)4
2,SSSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSSRqd='>Rj
',SSSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS;S2
SSSSMSC8CRoMNCs0HCRV;_d
SSSSVSH_Rc:H5VR5oEHE8N8sF-L0l0FDCHMR4<RnN2RM58RNs88I0H8E=R>R2c2RMoCC0sNCS
SSSSSNs00H0LkChRQQFaRVmR)vR c:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSSoLCHSM
SSSSSv)m :cRRv)m44nX
SSSSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSSRq.=q>R757).
2,SSSSSSSSSqSSd>R=R7q7)25d,S
SSSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSS2S;
SSSSCRM8oCCMsCN0R_HVcS;
SCSSMo8RCsMCNR0CLS;
SMSC8CRoMNCs0HCRV8_N8HsI8;0E
CSSMo8RCsMCNR0CH4V_n
8;S8CMRMoCC0sNCVRH_#d.;S

LR4:VRFsIMRHR04RFER5HdoE.MpHCRR-L0F0F.ldpCHM-2d./Rd.oCCMsCN0
LSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSNs00H0LkChRQQFaRVmR)vR 6:NRDLRCDHV#RkPMONID5*+d.L0F0F.ldpCHM,FRDI8N8sE,RHNoE8,8sR0LH,.Rd2S;
SHS#oDMNRbbHCF_8kR0#:0R#8F_Do;HO
LSSCMoH
SSS) mv6RR:)dmv.
X4SSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSq=4R>7Rq74)52S,
SSSSSqSS.>R=R7q7)25.,S
SSSSSSdSqRR=>q)775,d2
SSSSSSSSRqc=q>R757)c
2,SSSSSSSSm=RR>mR1zIa52H5L0S2
SSSSS;S2
CSSMo8RCsMCNR0CLS;
CRM8oCCMsCN0R;L4
H
SVn_4FH:RV5R5EEHodH.pM=CRRHREoHEpMRC2NRM85oEHEpd.HRMC>FRL0l0FdH.pM2C2RMoCC0sNCS
SLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SSo#HMRNDF_k0CRM8:0R#8F_Do;HO
SSSNs00H0LkChRQQFaRVmR)vR c:NRDLRCDHV#RkPMONED5HAoEFCs8s6-4,HREoFEAss8C-,46RoEHE8N8sL,RHR0,4;n2
LSSCMoH
SSS) mvcRR:)4mvn
X4SSSSSsbF0NRlbRR5qRjR=q>R757)j
2,SSSSSSSSq=4R>7Rq74)52S,
SSSSSqSS.>R=R7q7)25.,S
SSSSSSdSqRR=>q)775,d2
SSSSSSSSRmR=1>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./+d.4L25H
02SSSSS2SS;S
SCRM8oCCMsCN0R
L;S8CMRMoCC0sNCVRH_F4n;H
SVn_4#H:RV5R5EEHodH.pM<CRRHREoHEpMRC2NRM85oEHEpd.HRMC>FRL0l0FdH.pM2C2RMoCC0sNCS
SLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SSo#HMRNDF_k0CRM8:0R#8F_Do;HO
SSSNs00H0LkChRQQFaRVmR)vR 6:NRDLRCDHV#RkPMONED5HAoEFCs8s4-d,HREoFEAss8C-,d4RoEHE8N8sL,RHR0,d;.2
LSSCMoH
SSS) mv6RR:)dmv.
X4SSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSq=4R>7Rq74)52S,
SSSSSqSS.>R=R7q7)25.,S
SSSSSSdSqRR=>q)775,d2
SSSSSSSSRqc=q>R757)c
2,SSSSSSSSm=RR>mR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.50LH2S
SSSSSS
2;SMSC8CRoMNCs0LCR;C
SMo8RCsMCNR0CH4V_n
#;
RRRR_HVI0H8EH:RV0R5s0H#N_0CHRR<6o2RCsMCN
0CRRRRRRRRHFV_k:0jRRHV5oEHEpd.HRMC=FRL0l0FdH.pMRC2oCCMsCN0
RRRRRRRRRRRpamz5Rj2<1=Rm5zaj
2;RRRRRRRRCRM8oCCMsCN0R_HVFjk0;R
RRRRRRVRH_0Fk4H:RVER5HdoE.MpHCRR>L0F0F.ldpCHM2CRoMNCs0RC
RRRRRRRRRVRH_#ONCR4:H5VRL0F0FHlpM=CRR0LF0dFl.MpHCo2RCsMCN
0C-S-S#MHoN8DRHRVV:0R#8F_Do;HO
RSRRoLCH-M
-RRRRRRRRRRRR8RRHRVV<'=RjI'RERCMq)77RR<=Bemh_71a_tpmQeB_ mBa)45d+0LF0pFlH,MCR8N8s8IH0RE2
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#R''4;-
-SRRRRVRRFIs_HE80:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
S--RRRRRRRRRGlk0CsCRv:RznXw
S--SFSbsl0RN5bR
S--SRSSRRmR=p>Rm5zajH252-,
-SSSSQRRj>R=Rz1ma25j5,H2
S--SRSSRRQ4=1>Rm5za4H252-,
-SSSS1RRR>R=RV8HV-
-S2SS;-
-RRRRRRRRRRRRRMRC8CRoMNCs0VCRFIs_HE80;R
RRRRRRRRRRRRRpamz5Rj2<1=Rm5zajI2RERCMq)77RR<=Bemh_71a_tpmQeB_ mBa)45d+0LF0pFlH,MCR8N8s8IH0RE2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#1CRm5za4
2;RRRRRRRRRCRRMo8RCsMCNR0CHOV_N4#C;R
RRRRRRRRRR_HVOCN#.H:RVLR5FF00lMpHCRR>L0F0F.ldpCHM2CRoMNCs0-C
-#SSHNoMDHR8VRVj:0R#8F_Do;HO
RSRRCRLo
HM-R-RRRRRRRRRRRRR8VHVj=R<R''jRCIEM7Rq7<)R=mRBh1e_ap7_mBtQ_Be a5m)4L6+FF00lMpHCN,R8I8sHE802-R
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDC4R''-;
-RSRRRRRV_FsI0H8ERj:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0-C
-RSRRRRRRlRRksG0C:CRRXvzw-n
-SSSb0FsRblNR-5
-SSSSmRRR>R=Rzpma25j5,H2
S--SRSSRRQj=1>Rm5zajH252-,
-SSSSQRR4>R=Rz1ma2545,H2
S--SRSSRR1R=8>RHjVV
S--S;S2
R--RRRRRRRRRRRRR8CMRMoCC0sNCFRVsH_I8j0E;R
RRRRRRRRRRRRRpamz5Rj2<1=Rm5zajI2RERCMq)77RR<=Bemh_71a_tpmQeB_ mBa)654+0LF0pFlH,MCR8N8s8IH0RE2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#1CRm5za4
2;RRRRRRRRRCRRMo8RCsMCNR0CHOV_N.#C;R
RRRRRRMRC8CRoMNCs0HCRVk_F0
4;RRRRRRRRNV:RFIsRRRHM4FR0RH5Eo.EdpCHMRL-RFF00lpd.H-MCd/.2d4.-RMoCC0sNC-
-SHS#oDMNRV8HV:4RR8#0_oDFHPO_CFO0sE55HdoE.MpHCRR-L0F0F.ldpCHM-2d./-d.4FR8IFM0R;42
RSRRCRLo
HM-R-RRRRRRRRRRRRR8VHV425IRR<='Rj'IMECR7q7)RR<Bemh_71a_tpmQeB_ mBa).5d*+5I4L2+FF00lpd.H,MCR8N8s8IH0
E2-R-RRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C';4'
S--RRRRRFRVsH_I840E:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
S--RRRRRRRRRGlk0CsCRv:RznXw
S--SFSbsl0RN5bR
S--SRSSRRmR=p>Rm5zaIH252-,
-SSSSQRRj>R=Rzpma-5I4H252-,
-SSSSQRR4>R=Rz1ma+5I4H252-,
-SSSS1RRR>R=RV8HVI452-
-S2SS;-
-RRRRRRRRRRRRRMRC8CRoMNCs0VCRFIs_HE804R;
RRRRRRRRRRRRRzpma25IRR<=pamz54I-2ERICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)d5.*I2+4+0LF0dFl.MpHCN,R8I8sHE802R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C1amz54I+2R;
RRRRRCRRMo8RCsMCNR0CNR;
RRRRRR
RRRRRRVRH_#DN0:4nRRHV5H5Eo.EdpCHMRE=RHpoEH2MCR8NMRH5Eo.EdpCHMRL-RFF00lpd.HRMC>dRn2o2RCsMCN
0C-S-S#MHoN8DRH.VVR#:R0D8_FOoH;R
SRLRRCMoH
R--RRRRRRRRRRRRRV8HV<.R=jR''ERICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsC4s-6N,R8I8sHE802-R
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#'CR4
';-R-SRRRRRsVF_8IH0:E.RsVFRHHRMRRj0IFRHE80-o4RCsMCN
0C-R-SRRRRRRRRl0kGsRCC:zRvX
wn-S-SSsbF0NRlb
R5-S-SSRSRm=RR>mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d5.2H
2,-S-SSRSRQ=jR>mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d4.-225H,-
-SSSSR4RQRR=>1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.H252-,
-SSSS1RRR>R=RV8HV-.
-SSS2-;
-RRRRRRRRRRRRCRRMo8RCsMCNR0CV_FsI0H8E
.;RRRRRRRRRRRRpamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d2=R<RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.2-4RS
SSISSERCMq)77RB<Rm_he1_a7pQmtB _eB)am5oEHEsAF8-Cs4R6,Ns88I0H8ER2
RRRRRRRRRRRRRRRRRCRRDR#C1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.
2;RRRRRRRRCRM8oCCMsCN0R_HVD0N#4
n;
RRRRRRRR_HVD0N#dR.:H5VR5oEHEpd.HRMC<ERRHpoEH2MCR8NMRH5Eo.EdpCHMRL-RFF00lpd.HRMC>dRn2o2RCsMCN
0C-S-S#MHoN8DRHdVVR#:R0D8_FOoH;R
SRLRRCMoH
R--RRRRRRRRRRRRRV8HV<dR=jR''ERICqMR7R7)<mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCds-4N,R8I8sHE802-R
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#'CR4
';-R-SRRRRRsVF_8IH0:EdRsVFRHHRMRRj0IFRHE80-o4RCsMCN
0C-R-SRRRRRRRRl0kGsRCC:zRvX
wn-S-SSsbF0NRlb
R5-S-SSRSRm=RR>mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d5.2H
2,-S-SSRSRQ=jR>mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d4.-225H,-
-SSSSR4RQRR=>1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.H252-,
-SSSS1RRR>R=RV8HV-d
-SSS2-;
-RRRRRRRRRRRRCRRMo8RCsMCNR0CV_FsI0H8E
d;RRRRRRRRRRRRpamz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d2=R<RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.2-4RS
SSISSERCMq)77RB<Rm_he1_a7pQmtB _eB)am5oEHEsAF8-CsdR4,Ns88I0H8ER2
RRRRRRRRRRRRRRRRRCRRDR#C1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.
2;RRRRRRRRCRM8oCCMsCN0R_HVD0N#d
.;
RRRRRRRR_HVF.k0:VRHRH5EoFEAss8CRL-RFF00lMpHCRR<nRc2oCCMsCN0
RRRRRRRRRRRR7RRm_zaNRkG<8=RVRD0IMECRR5RRqR57R7)>mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFs57q7)RR<Bemh_71a_tpmQeB_ mBa)F5L0l0FpCHM,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#pCRm5zaj
2;RRRRRRRRCRM8oCCMsCN0R_HVF.k0;R
RRRRRRVRH_0FkdH:RVER5HAoEFCs8sRR-L0F0FHlpM>CRR2ndRMoCC0sNCR
RRRRRRRRRRRRR7amz_GNkRR<=80VDRCIEMRR5R5RRq)77RB>Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRRsqR57R7)<mRBh1e_ap7_mBtQ_Be a5m)L0F0FHlpMRC,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.
2;RRRRRRRRCRM8oCCMsCN0R_HVFdk0;R
RRCRRMo8RCsMCNR0CHIV_HE80;R
RRR
RRHRRVH_I8j0E:VRHRs50HN#00HC_RR>=6o2RCsMCN
0CRRRRRRRRHOV_N4#C:VRHRF5L0l0FpCHMRL=RFF00lpd.H2MCRMoCC0sNCR
RRRRRRRRRRz7mak_NG=R<Rz1ma25jRCIEMRR5R5RRq)77RR<=Bemh_71a_tpmQeB_ mBa)45d+0LF0pFlH,MCR8N8s8IH02E2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRM58Rq)77RR>=Bemh_71a_tpmQeB_ mBa)F5L0l0FpCHM,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CHOV_N4#C;R
RRRRRRVRH_#ONCR.:H5VRL0F0FHlpM>CRR0LF0dFl.MpHCo2RCsMCN
0CRRRRRRRRR7RRm_zaNRkG<1=Rm5zajI2RERCM5RRRR75q7<)R=mRBh1e_ap7_mBtQ_Be a5m)4L6+FF00lMpHCN,R8I8sHE802
2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNSRM58Rq)77RR>=Bemh_71a_tpmQeB_ mBa)F5L0l0FpCHM,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CHOV_N.#C;R
RRRRRRjRN:FRVsRRIH4MRRR0F5oEHEpd.H-MCL0F0F.ldpCHM-2d./Rd.oCCMsCN0
RRRRRRRRRRRR7RRm_zaNRkG<1=Rm5zaII2RERCM5RRRR75q7<)R=mRBh1e_ap7_mBtQ_Be a5m)d5.*I2+4+FRL0l0FdH.pM4C-,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN8qR57R7)>B=Rm_he1_a7pQmtB _eB)am5*d.IF+L0l0FdH.pMRC,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R;Nj
RRRRRRRR_HV#dkb.H:RV5R5EEHodH.pM=CRRHREoHEpMRC2NRM85oEHEpd.HRMC-FRL0l0FdH.pM>CRR2nd2CRoMNCs0RC
RRRRRRRRRRRRRz7mak_NG=R<Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2dR.2
SSSRSRSSESIC5MRRRRR57q7)=R<RhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8NMR75q7>)R=mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsC4s-6N,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_b#kd
.;RRRRRRRRH#V_knb4:VRHRE55HdoE.MpHCRR<RoEHEMpHCN2RM58REEHodH.pM-CRR0LF0dFl.MpHCRR>n2d2RMoCC0sNCR
RRRRRRRRRRRRR7amz_GNkRR<=1amz5H5Eo.EdpCHM-0LF0dFl.MpHCd2/.
2RSRSSRSSSSCIEMRR5R5RRq)77RR<=Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRM857q7)=R>RhBmea_17m_pt_QBea BmE)5HAoEFCs8s4-d,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HV#4kbnR;
RRRRRHRRVF_DIH:RVLR5FF00lMpHCRR>jo2RCsMCN
0CRRRRRRRRR7RRm_zaNRkG<8=RVRD0IMECRR5RR75q7<)RRhBmea_17m_pt_QBea BmL)5FF00lMpHCN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSRF5sRq)77RB>Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CHDV_F
I;RRRRRRRRHDV_F:IjRRHV50LF0pFlHRMC<2R4RMoCC0sNCR
RRRRRRRRRRz7mak_NG=R<RD8V0ERIC5MRq)77RB>Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVF_DI
j;RRRRR8CMRMoCC0sNCVRH_8IH0;Ej
M
C8sRNO0EHCkO0s#CRCODC0m_)v
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCFRIso	3CNMbOo	NCD3ND
;
DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$)RmvHS#
oCCMsRHO5S
SSlVNHRD$:0R#soHMRR:="$NM"S;
SHSI8R0E:MRH0CCos=R:R
c;SNSS8I8sHE80RH:RMo0CC:sR=;R(
SSSDNFI8R8s:MRH0CCos=R:R
j;SESSHNoE8R8s:MRH0CCos=R:R;(U
SSS0DNLCRR:s0FlNCLD;S
SSD8V0RR:sIFlF
s8S
2;SsbF0
R5SqSS7R7):MRHR8#0_oDFHPO_CFO0sNR58I8sHE80R4-RRI8FMR0Fj
2;S7SSmRza:kRF00R#8F_Do_HOP0COF5sRI0H8ERR-4FR8IFM0R
j2S;S2
N
S0H0sLCk0Rs\3N\M	RH:RMo0CC
s;RRRRNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MC8RM00H$mR)v
;
NEsOHO0C0CksRD#CC_O0)RmvF)VRmHvR#O
SFFlbM0CMRv)m_#LNCS
SoCCMsRHO5S
SSHSI8R0E:MRH0CCosS;
SNSS8I8sHE80RH:RMo0CC
s;SSSSDNFI8R8s:MRH0CCosS;
SESSHNoE8R8s:MRH0CCosS;
S0SSNCLDRs:RFNl0L;DC
SSSSD8V0RR:sIFlF
s8S;S2
bSSFRs05S
SS7Sq7:)RRRHM#_08DHFoOC_POs0FR85N8HsI8R0E-RR48MFI0jFR2S;
S7SSmRza:kRF00R#8F_Do_HOP0COF5sRI0H8ERR-4FR8IFM0R
j2S2SS;C
SMO8RFFlbM0CM;S

O#FM00NMRLM0RH:RMo0CC:sR=nR4;S

VOkM0MHFRN#0sF0)lMpHCCRs0MksR0HMCsoCR
H#SNSPsLHND#CRHRxC:MRH0CCosS;
SMOF#M0N0DRLF#O	HRxC:MRH0CCos=R:RLM0Rn*RcS;
LHCoMS
SH5VRDNFI8R8slRF8LODF	x#HC=2RRRRj0MEC
SSSskC0sDMRF8IN8+sRRFLDOH	#x
C;SDSC#SC
SCSs0MksRD55F8IN8+sRRFLDOH	#x-CRRR42/DRLF#O	H2xCRL*RD	FO#CHx;S
SCRM8H
V;S8CMRMVkOF0HM0R#N)s0FHlpM
C;
FSOMN#0ML0RD	FO#CHxRH:RMo0CC:sR=cRnRM*R0
L;SMOF#M0N0HRDl8q8sRR:HCM0oRCs:#=R00Ns)pFlH;MCRO
SF0M#NRM0MsL_FVl_sRNO:MRH0CCos=R:RH5Eo8EN8-sRRlDHqs88R4+R2L/RD	FO#CHx;O
SF0M#NRM0D0CV_lsF_NVsORR:HCM0oRCs:5=REEHoNs88RD-RH8lq8+sRRR42lRF8LODF	x#HC
;
Sb0$CNR0L_DC80FkRRH#NNss$MR5LF_sls_VN4O+RI8FMR0FjF2RVFRslsIF8
;
So#HMRND80Fk_lsFR0:RNCLD_k8F0L;
CMoH
H
SVH_Lov)m:VRHRH5Eo8EN8-sRRIDFNs88R4+RRL>RD	FO#CHx2CRoMNCs0SC
So#HMRND80Fk_sVH#R0,7amz_GNkRs:RFFlIs
8;SHS#oDMNR7q7)k_NGq,R7_7)VRR:#_08DHFoOC_POs0FR85N8HsI8R0E-RR48MFI0jFR2S;
LHCoMS

SsVF_bbHCV:RFHsRRRHMjFR0R8N8s8IH04E-RMoCC0sNCS
SS0N0skHL0\CR3MsN	F\RVCRsoR#q:NRDLRCDHj#R;S
SS0N0skHL0\CR3MsN	F\RVCRsoR#A:NRDLRCDH4#R;R
RRRRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:qRRLDNCHDR#;R4
RRRRRRRRRRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoARR:DCNLD#RHR
4;SCSLo
HMSsSSCqo#:HRbbkCLVS
SSsbF0NRlbS5
SSSSR=QR>7Rq7H)52S,
SRSSSRRm=q>R7_7)V25H
SSSS;S2
S
SSosC#RA:bCHbL
kVSbSSFRs0l5Nb
SSSSQSRRR=>q)77_HV52S,
SRSSSRRm=q>R7_7)N5kGHS2
SSSS2S;
S8CMRMoCC0sNCFRVsH_bb
C;
)SSm4v (RR:)_mvLCN#
SSSoCCMsRHOl5Nb
SSSS8IH0SERSR=>I0H8ES,
SNSS8I8sHE80R=RS>8RN8HsI8,0ERS
SSFSDI8N8sRRRSR=>DNFI8,8s
SSSSoEHE8N8sRRRSR=>DqHl8-8s4S,
S0SSNCLDRSRR=0>RNCLD,S
SSVS8DR0RR=SS>VR8DS0
S
S2SbSSFRs0lRNb5qRR7R7)=q>R7_7)V
,RSSSSSmS7z=aR>FR8kV0_H0s#
SSSS;S2SS

Sk8F0F_sl25jRR<=80Fk_sVH#I0RERCM57q7)k_NG=R>RhBmea_17m_pt_QBea BmD)5F8IN8Rs,Ns88I0H8E
22SSSSSSSSRCRRDR#C80VD;S

SsVF_FDFbV:RFHsRRRHM4FR0R_MLs_FlVOsNRMoCC0sNCS
SSo#HMRND80Fk_N#0o:CRRlsFI8Fs;S
SLHCoMS
SSv)m :6RRv)m_#LNCS
SSMoCCOsHRblN5S
SSHSI8R0ES>S=R8IH0
E,SSSSNs88I0H8ESRR=N>R8I8sHE80,SR
SDSSF8IN8RsRR>S=RlDHqs88R5+RH2-4*FLDOH	#x
C,SSSSEEHoNs88RSRR=D>RH8lq8+sRRLH*D	FO#CHx-R4,
SSSSL0NDRCRR>S=RL0ND
C,SSSS80VDRSRRSR=>80VD
SSS2S
SSsbF0NRlbRR5R7q7)>R=R7q7),_VRS
SSSSS7amzRR=>80Fk_N#0oSC
SSSS2
;S
SSS80Fk_lsF5RH2<8=RF_k0#o0NCERIC5MRq)77_GNkRR>=Bemh_71a_tpmQeB_ mBa)H5Dl8q8sH+5-*42LODF	x#HCN,R8I8sHE802S2
SSSSSRSSRDRC#8CRF_k0s5FlH2-4;S
SCRM8oCCMsCN0RsVF_FDFbS;

HSSVH_#xRC:H5VRD0CV_lsF_NVsORR>jo2RCsMCN
0CS#SSHNoMDFR8k#0_0CNoRs:RFFlIs
8;SCSLo
HMS)SSm6v R):RmLv_N
#CSoSSCsMCHlORN
b5SSSSI0H8ESRS=I>RHE80,S
SS8SN8HsI8R0ER>S=R8N8s8IH0RE,
SSSSIDFNs88RSRR=D>RH8lq8+sRR_MLs_FlVOsN*FLDOH	#x
C,SSSSEEHoNs88RSRR=E>RHNoE8,8sRS
SSNS0LRDCR=RS>NR0L,DC
SSSSD8V0RRRS>S=RD8V0S
SSS2
SFSbsl0RN5bRR7Rq7=)R>7Rq7V)_,SR
SSSSSz7ma>R=Rk8F00_#N
oCSSSSSS2;
SS
SFS8ks0_FMl5LF_sls_VN4O+2=R<Rk8F0F_slL5M_lsF_NVsOS2
SSSSSSSSSESIC5MRq)77_GNkRB<Rm_he1_a7pQmtB _eB)am5lDHqs88+_MLs_FlVOsN*FLDOH	#xRC,Ns88I0H8E
22SSSSSSSSRSRRSRRRR#CDCFR8k#0_0CNo;

SS7SSm_zaNRkG<8=RVRD0IMECR75q7N)_k>GRRhBmea_17m_pt_QBea BmE)5HNoE8,8sR8N8s8IH02E2
SSSSSSSR#CDCFR8ks0_FMl5LF_sls_VN4O+2S;
S8CMRMoCC0sNCVRH_x#HCS;

HSSV#_MH:xCRRHV5VDC0F_sls_VN=ORRRj2oCCMsCN0
SSS7amz_GNkRR<=80VDRCIEMqR57_7)NRkG>mRBh1e_ap7_mBtQ_Be a5m)EEHoNs88,8RN8HsI820E2S
SSSSSSDRC#8CRF_k0s5FlMsL_FVl_s2NO;S
SCRM8oCCMsCN0R_HVMx#HC
;
SFSVsH_bbRC:VRFsHMRHR0jRFHRI8-0E4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRCRo#:NRDLRCDH.#R;R
RRRRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;SLSRCMoH
SSSRosC#b:RHLbCkSV
SRSSb0FsRblN5S
SRSRRSRSSR=QR>mR7zNa_kHG52S,
SRRRSSSSRRRm=7>Rm5zaHS2
SSSSS;R2
RSSCRM8oCCMsCN0RsVF_bbHC
;
S8CMRMoCC0sNCVRH_oLH);mv
H
SVl_#N)DDmRv:H5VREEHoNs88RD-RF8IN8+sRR<4R=DRLF#O	H2xCRMoCC0sNCS
S#MHoNqDR7_7)VRR:#_08DHFoOC_POs0FR85N8HsI8R0E-RR48MFI0jFR2S;
LHCoMS
SV_FsbCHb:FRVsRRHHjMRRR0FNs88I0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#CoqRR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:qRRLDNCHDR#;R4
LSSCMoH
SSSs#Coqb:RHLbCkSV
SbSSFRs0l5Nb
SSSSRSQ=q>R757)H
2,SSSSS=mR>7Rq7V)_5
H2SSSS2S;
S8CMRMoCC0sNCFRVsH_bb
C;
mS)vR 6:mR)vN_L#SC
SoSSCsMCHlORN
b5SSSSSISSHE80R=SS>HRI8,0E
SRRSSSSS8SN8HsI8R0ER>R=R8N8s8IH0RE,
SSSSSSSDNFI8R8sR=RS>FRDI8N8sS,
SSSSSHSEo8EN8RsRR>S=RoEHE8N8sS,
SSSSSNS0LRDCR=RS>NR0L,DC
SSSSSSS80VDRSRRSR=>80VD
SSSSSSS2S
SSFSbsl0RN5bRR7Rq7=)R>7Rq7V)_,SR
SSSSSmS7z=aR>mR7zSa
SSSSSS2;
C
SMo8RCsMCNR0CH#V_lDND);mv
M
C8sRNO0EHCkO0s#CRCODC0m_)v
;

