-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRRRR:RwCHG8FRuHRM0NRM8wNDF0oHMRHuFM00R$#bCRObN	CNo

---R-RRLpHs$NsR:RRRERaHb#RNNO	o#CREDNDRRLCObFlH8DCR0HMFRRNDsHLNRs$
R--RRRRRRRRRRRRR#RR$FlLDNHODRD$MCNl8 RQ R 3

---R-RRP7CCbDFC:s#RORqODCDCRsNep]7-RaBNRM8Q   Rju4(WnRFHs	MtoRsbFk

---R-RRsukbCF#R:RRRCR7VHHM0MHF#FRVs#RkCMRHRGVHCb8RF0HMR8NMRFVDNM0HoFRbH
M0-R-RRRRRRRRRRRRRRsRNHl0ECO0HRObN	CNo#-
-
R--RFRh0RCRRRRR:aRRERH#b	NONRoClRN$LlCRFV8HHRC80HFRMkOD8NCR808HHNFMDNR80-N
-RRRRRRRRRRRRRR:RJsCkCHs8$RLRF0FDR#,LRk0Hl0RkR#0HMMRFNRI$ERONCMoRC0E
R--RRRRRRRRRRRR:CRRGs0CMRNDHCM0sOVNCF#RsHR#lNkD0MHFRELCNFPHsVRFRC0E
R--RRRRRRRRRRRR:8RRCs#OHHb0FRM3QH0R#CRbs#lH#DHLCFR0R8N8RlOFl0CM#MRN8s/F
R--RRRRRRRRRRRR:NRR0H0sLCk0#FR0RC0ERObN	CNoRO8CDNNs0MHF#L,RkM0RF00RFERONCMo
R--RRRRRRRRRRRR:FRRsCR8DCC0R$NMRHFsoNHMDHRDMRC#F0VREbCRNNO	o8CRCNODsHN0F
M3-R-RRRRRRRRRR:RRRERaCNRbOo	NCFRL8l$RNL$RCERONCMo8MRFDH$RMORNO8FsNCMOR0IHE-
-RRRRRRRRRRRRRR:R0REC0lCs#VRFRNBDkR#C4FnRVER0H##R08NMN3s8
R--RRRRRRRRRRRR:-
-R---------------------------------------------------------------------
-RCf)PHH#FRM:4j..R-f
-7RfN:0CRj.jUc-j-R4j44(:ng:jRg+jd5jRa,EkRR4jqRbs.Ujj2
Rf---R-----------------------------------------------------------------
--
ObN	CNoRGVHCV8_D0FN_b0$CH#R#R

RR--aC$b##RkCV8RFosRCsMCHRO#FVVRH8GC_MoCCOsH_ob	

RRR$R0bVCRH8GC_ksFM#8_0C$D_b0$C#RHRH5VG_C8sMFk8V,RH8GC_k0sM0ONC
2;RRR
Rb0$CHRVG_C8FsPCVIDF_$#0D0C_$RbCH5#RVCHG8N_#0Nks0RC,VCHG8s_IN;b2
R
R-a-R$RbCk8#CRsVFRMoCCOsH#VRFRFVDNo0_CsMCHbO_	
o
R-R-RCaE#NCRs0CRE#CRNRlCN0#REBCRR_w a mhq1) aw,R u_zW7q), Rw_W7mh)Wq7R,
RR--NRM8wa _m)Wq7)Z mDRVFHN0MboRF0HMRksFMM8HoNRlO#sF3R

Rb0$CFRsk_M80C$bRRH#5ksFMM8_CCNs#R0,R-RR-CR7VDNk0M,RCCNs#p0R1'ARjR'
RRRRRRRRRRRRRRRRRRRRRksFMH8_MRV,RRRRR-RR-FR)kRM80NFIsb8RF0#HHRPCHHMVM$H0
RRRRRRRRRRRRRRRRRRRRsRRF8kM_oMCH,MVRRRRRR--)MFk8FR0I8NsRoMCNP0HCMRHVHHM0R$
RRRRRRRRRRRRRRRRRRRRRksFMx8_C2sF;RRRR-RR-FR)kRM80NFIsx8RCRsF5k0sM0ONC
2
CRM8b	NONRoCVCHG8D_VF_N00C$b#
;

