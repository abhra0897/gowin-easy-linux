`ifndef AE250_SMU_CONST_VH
`define AE250_SMU_CONST_VH

//`define AE250_SMU_RESET_VECTOR_DEFAULT	32'h8000_0000

`define AE250_SMU_CCLKE_DEFAULT		1'b1
`define AE250_SMU_HCLKE_DEFAULT		1'b1
`define AE250_SMU_PCLKE_DEFAULT		1'b1
`define AE250_SMU_CLKE_DEFAULT		{8'h00, `AE250_SMU_PCLKE_DEFAULT, `AE250_SMU_HCLKE_DEFAULT, `AE250_SMU_CCLKE_DEFAULT}

`ifdef AE250_CLK_RATIO_4_4_2
	`define AE250_SMU_CLKR_DEFAULT		4'h2
`elsif AE250_CLK_RATIO_4_4_1
	`define AE250_SMU_CLKR_DEFAULT		4'h4
`elsif AE250_CLK_RATIO_4_2_2
	`define AE250_SMU_CLKR_DEFAULT		4'h6
`elsif AE250_CLK_RATIO_4_2_1
	`define AE250_SMU_CLKR_DEFAULT		4'h8
`else
	`define AE250_SMU_CLKR_DEFAULT		4'h0
`endif


`endif
