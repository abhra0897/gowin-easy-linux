`ifndef ATCRTC100_CONST_VH
`define ATCRTC100_CONST_VH

`define ATCRTC100_PRODUCT_ID	32'h03011006

`ifdef ATCRTC100_HALF_SECOND_SUPPORT
	`define ATCRTC100_DIVIDER_WIDTH	14
	`define	ATCRTC100_SEC_WIDTH	7
	`define ATCRTC100_ST_WIDTH	8
`else
	`define ATCRTC100_DIVIDER_WIDTH	15
	`define ATCRTC100_SEC_WIDTH	6
	`define ATCRTC100_ST_WIDTH      7
`endif
`define ATCRTC100_CTL_WIDTH	9

`define ATCRTC100_SDO_SEC_WIDTH	6
`define	ATCRTC100_MIN_WIDTH	6
`define	ATCRTC100_HOUR_WIDTH	5
`define	ATCRTC100_DAY_WIDTH	`ATCRTC100_DAY_BITS

`define ATCRTC100_SDO_WIDTH 	(`ATCRTC100_SDO_SEC_WIDTH + `ATCRTC100_MIN_WIDTH + `ATCRTC100_HOUR_WIDTH + `ATCRTC100_DAY_WIDTH)
`define ATCRTC100_ALM_WIDTH	(`ATCRTC100_SDO_SEC_WIDTH + `ATCRTC100_MIN_WIDTH + `ATCRTC100_HOUR_WIDTH)

`endif
