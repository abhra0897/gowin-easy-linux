//------------------------------------------------------------------------
// Filename     : atcapbbrg100_config.vh
// Description  : specify APB bridge configurations
//------------------------------------------------------------------------
`ifndef ATCAPBBRG100_CONFIG
`define ATCAPBBRG100_CONFIG

// Specify APB slaves according to SoC configuration
`include "ae250_config.vh"
`include "ae250_const.vh"

`define ATCAPBBRG100_SLV_1

`ifdef AE250_UART1_SUPPORT
	`define	ATCAPBBRG100_SLV_2
`endif

`ifdef AE250_UART2_SUPPORT
	`define	ATCAPBBRG100_SLV_3
`endif

`ifdef AE250_PIT_SUPPORT
	`define ATCAPBBRG100_SLV_4
`endif

`ifdef AE250_WDT_SUPPORT
	`define ATCAPBBRG100_SLV_5
`endif

`ifdef AE250_RTC_SUPPORT
`define ATCAPBBRG100_SLV_6
`endif

`ifdef AE250_GPIO_SUPPORT
`define ATCAPBBRG100_SLV_7
`endif

`ifdef AE250_I2C_SUPPORT
	`define	ATCAPBBRG100_SLV_8
`endif

`ifdef AE250_SPI1_SUPPORT
	`define	ATCAPBBRG100_SLV_9
`endif

`ifdef AE250_SPI2_SUPPORT
	`define	ATCAPBBRG100_SLV_10
`endif

`ifdef AE250_SDC_SUPPORT
	`define	ATCAPBBRG100_SLV_11
`endif

`ifdef AE250_SPI3_SUPPORT
	`define	ATCAPBBRG100_SLV_13
`endif

`ifdef AE250_SPI4_SUPPORT
	`define	ATCAPBBRG100_SLV_14
`endif

`ifdef AE250_I2C2_SUPPORT	// For CF1
	`define	ATCAPBBRG100_SLV_16
`endif

`ifdef AE250_PIT2_SUPPORT	// For CF1
	`define	ATCAPBBRG100_SLV_17
`endif

`ifdef AE250_PIT3_SUPPORT	// For CF1
	`define	ATCAPBBRG100_SLV_18
`endif

`ifdef AE250_PIT4_SUPPORT	// For CF1
	`define	ATCAPBBRG100_SLV_19
`endif

`ifdef AE250_PIT5_SUPPORT	// For CF1
	`define	ATCAPBBRG100_SLV_20
`endif


`ifdef ATCAPBBRG100_ADDR_WIDTH_24
	`define	ATCAPBBRG100_ADDR_DECODE_WIDTH	17
	`define	ATCAPBBRG100_SLV1_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h01000
	`define	ATCAPBBRG100_SLV2_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h02000
	`define	ATCAPBBRG100_SLV3_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h03000
	`define	ATCAPBBRG100_SLV4_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h04000
	`define	ATCAPBBRG100_SLV5_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h05000
	`define	ATCAPBBRG100_SLV6_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h06000
	`define	ATCAPBBRG100_SLV7_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h07000
	`define	ATCAPBBRG100_SLV8_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0a000
	`define	ATCAPBBRG100_SLV9_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0b000
	`define	ATCAPBBRG100_SLV10_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0f000
	`define	ATCAPBBRG100_SLV11_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0e000
	`define	ATCAPBBRG100_SLV12_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h11000

	// CF1
	`define	ATCAPBBRG100_SLV13_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h19000
	`define	ATCAPBBRG100_SLV14_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1a000
	`define	ATCAPBBRG100_SLV16_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1b000
	`define	ATCAPBBRG100_SLV17_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h10000
	`define	ATCAPBBRG100_SLV18_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h11000
	`define	ATCAPBBRG100_SLV19_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h12000
	`define	ATCAPBBRG100_SLV20_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h13000

	`define	ATCAPBBRG100_SLV1_SIZE		3
	`define	ATCAPBBRG100_SLV2_SIZE		3
	`define	ATCAPBBRG100_SLV3_SIZE		3
	`define	ATCAPBBRG100_SLV4_SIZE		3
	`define	ATCAPBBRG100_SLV5_SIZE		3
	`define	ATCAPBBRG100_SLV6_SIZE		3
	`define	ATCAPBBRG100_SLV7_SIZE		3
	`define	ATCAPBBRG100_SLV8_SIZE		3
	`define	ATCAPBBRG100_SLV9_SIZE		3
	`define	ATCAPBBRG100_SLV10_SIZE		3
	`define	ATCAPBBRG100_SLV11_SIZE		3
	`define	ATCAPBBRG100_SLV12_SIZE		3

	// CF1
	`define	ATCAPBBRG100_SLV13_SIZE		3
	`define	ATCAPBBRG100_SLV14_SIZE		3
	`define	ATCAPBBRG100_SLV16_SIZE		3
	`define	ATCAPBBRG100_SLV17_SIZE		3
	`define	ATCAPBBRG100_SLV18_SIZE		3
	`define	ATCAPBBRG100_SLV19_SIZE		3
	`define	ATCAPBBRG100_SLV20_SIZE		3
`else	// !ATCAPBBRG100_ADDR_WIDTH_24
	`define	ATCAPBBRG100_ADDR_DECODE_WIDTH	25
	//`define	ATCAPBBRG100_SLV1_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0100000	// SMU
	//`define	ATCAPBBRG100_SLV2_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0200000	// UART1
	//`define	ATCAPBBRG100_SLV3_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0300000	// UART2
	//`define	ATCAPBBRG100_SLV4_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0400000	// PIT
	//`define	ATCAPBBRG100_SLV5_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0500000	// WDT
	//`define	ATCAPBBRG100_SLV6_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0600000	// RTC
	//`define	ATCAPBBRG100_SLV7_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0700000	// GPIO
	//`define	ATCAPBBRG100_SLV8_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0a00000	// I2C
	//`define	ATCAPBBRG100_SLV9_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0b00000	// SPI1
	//`define	ATCAPBBRG100_SLV10_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0f00000	// SPI2
	`define	ATCAPBBRG100_SLV11_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0e00000	// SDC
	`define	ATCAPBBRG100_SLV12_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1100000	// Unused now

	// CF1
	`define	ATCAPBBRG100_SLV13_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1900000	// SPI3
	`define	ATCAPBBRG100_SLV14_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1a00000	// SPI4
	`define	ATCAPBBRG100_SLV16_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1b00000	// I2C2
	`define	ATCAPBBRG100_SLV17_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1000000	// PIT2
	`define	ATCAPBBRG100_SLV18_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1100000	// PIT3
	`define	ATCAPBBRG100_SLV19_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1200000	// PIT4
	`define	ATCAPBBRG100_SLV20_OFFSET	`ATCAPBBRG100_ADDR_DECODE_WIDTH'h1300000	// PIT5

	`define	ATCAPBBRG100_SLV1_SIZE		1
	`define	ATCAPBBRG100_SLV2_SIZE		1
	`define	ATCAPBBRG100_SLV3_SIZE		1
	`define	ATCAPBBRG100_SLV4_SIZE		1
	`define	ATCAPBBRG100_SLV5_SIZE		1
	`define	ATCAPBBRG100_SLV6_SIZE		1
	`define	ATCAPBBRG100_SLV7_SIZE		1
	`define	ATCAPBBRG100_SLV8_SIZE		1
	`define	ATCAPBBRG100_SLV9_SIZE		1
	`define	ATCAPBBRG100_SLV10_SIZE		1
	`define	ATCAPBBRG100_SLV11_SIZE		1
	`define	ATCAPBBRG100_SLV12_SIZE		1

	// CF1
	`define	ATCAPBBRG100_SLV13_SIZE		1
	`define	ATCAPBBRG100_SLV14_SIZE		1
	`define	ATCAPBBRG100_SLV16_SIZE		1
	`define	ATCAPBBRG100_SLV17_SIZE		1
	`define	ATCAPBBRG100_SLV18_SIZE		1
	`define	ATCAPBBRG100_SLV19_SIZE		1
	`define	ATCAPBBRG100_SLV20_SIZE		1
`endif	// !ATCAPBBRG100_ADDR_WIDTH_24

`endif	// !ATCAPBBRG100_CONFIG
