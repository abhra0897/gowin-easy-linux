@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ha_ "Xa;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"
`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vtR

RHHM0DHNRoLCHRM
RHRRVMR5kOl_	<#R=2RjRoLCHRM
RRRRRDFP_sCsF0s_5D"QDNCoDNRPDRkCVRFsbNNslCC0skRMl	_O#ERIHROEl0k#RRLC#RC00PFRNCDkRCosNs0CRN0EM"Rj2R;
RCRRMR8
R8CM
H
`VV8CRpme_q1])_ 7B m7
R
RHCM0oRCsHRR=j
;
RDRNI#N$RR@@5#bFCC8oR	OD2CRLo
HMRRRRH5VR`pme_1)  1a_Qqthp=R!RL4'jL2RCMoH
RRRRHRRV#R500Ns_CCPM=0R='R4LR42LHCoMR
RRRRRRRRH<M=RkOl_	
#;RRRRRMRC8RR
RRRRR#CDCVRHRR5H>2R4RoLCHRM
RRRRRHRRRR<=HRR-4R;
RRRRR8CM
RRRR8CM
RRRR#CDCCRLo
HMRRRRRRRH<j=R;R
RRMRC8R
RC
M8
M`C8RHV/m/Re1p_] q)7m_B7
 
`8HVCmVReqp_1)1 ah_m
R
RbbsFC$s0R1q1 _)aha X_q1a)Wa_Qma]zaa_ _1auR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RN#0sC0_P0CMR>|-RMyykOl_	0#RC_#0CsGb;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)ha_ _Xaaa 1_aWQ]amz_q1a)ua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RMRF05#5!00Ns_CCPMR02ykyMl	_O#CR0#C0_G2bs;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)ha_ _Xahmm_ep )quu_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R#s0N0P_CCRM0|R->5<HR=2R4;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_Xh aZ_X__mh1)aqae_  _hauR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R55!fkH#MF	MI#M500Ns_CCPM2022R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aha X__XZmah_ _1a )Xu_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42ROR5E	CO_#lH#oHM_N#0s|0R|bRfN5#0#s0N0P_CC,M0M_klO2	#2-R|>!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRM_klOR	#>2RjRoLCH:MRRNN_#s#C0C_MG#0_00Ns_0IHE0Fk_#0C0R
RRRRRRRRRq1_q1a )_Xh aa_1q_)aW]Qam_zaaa 1_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _hX1a_aaq)_aWQ]amz_1a a2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRRH#MRF0NC##s80CR0NVCCsRD#NbCVRFRlMk_#O	ROO$DRC#VlsFRN#0sC0RP0CM"
2;
RRRRRRRRHRRVOR5E	CO_#lH#oHM_N#0sR02LHCoMRR:N#_N#0Cs_GMC0C_0#I0_HF0Ek#0_00Ns
RRRRRRRRRRRRqq_1)1 a _hXaa_ _1aW]Qam_za1)aqa:_u
RRRRRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Xh a _a1Wa_Qma]z1a_aaq)_
u2RRRRRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#M#FRRH#NC##s80CRHRI0kEF0RRNOsFsCF#bMM8Ho0R#N_s0CMPC0;"2
RRRRRRRRCRRMR8
RRRRRRRRRRHV5E!OC_O	FsPCDbNbH2MoRoLCH:MRRNN_#s#C0C_MGM0_FP_FCNsDbR
RRRRRRRRRR_Rqq 11)ha_ _Xahmm_ep )quu_:R
RRRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _hXha_me_m q)pu2_u
RRRRRRRRRRRR#CDCPRFDs_Cs_Fs0Q5"DoDCNFDRPDCsNHbbMOoRFHM80MHFRRFV#s0N0PRCCRM0H8#RCO0C0"C82R;
RRRRRRRRR8CM
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRR_Rqq 11)ha_ _XaXmZ_ha_1q_)a he a:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)ha_ _XaXmZ_ha_1q_)a he a2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N#0sC0_P0CMRMOF0MNH#RRXFZsR"
2;
RRRRRRRRqRR_1q1 _)aha X__XZmah_ _1a )Xu_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _hXXa_Zh_m_1a aX_ uu)_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRC
M8RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRRHV5lMk_#O	Rj>R2CRLoRHM:_RlNC##sM0_C_G0#s0N0H_I0kEF0C_0#R0
RRRRRRRRRqv_1)1 a _hX1a_aaq)_aWQ]amz_1a a:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)ha_ _Xa1)aqaQ_Waz]ma _a1ua_2
;
RRRRRRRRRVRHRE5OC_O	l#H#H_Mo#s0N0L2RCMoHRl:R_#N#C_s0M0CG_#0C0H_I0kEF00_#N
s0RRRRRRRRRRRRv1_q1a )_Xh a _a1Wa_Qma]z1a_aaq)_
u:RRRRRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aha X_1a aQ_Waz]maa_1q_)au
2;RRRRRRRRRMRC8R
RRRRRRRRRH5VR!COEOF	_PDCsNHbbMRo2LHCoMRR:l#_N#0Cs_GMC0F_M_CFPsbDN
RRRRRRRRRRRRqv_1)1 a _hXha_me_m q)pu:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Xh am_h_ me)upq_;u2
RRRRRRRRCRRM
8

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRRRRRv1_q1a )_Xh aZ_X__mh1)aqae_  _hauR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Xh aZ_X__mh1)aqae_  _hau
2;
RRRRRRRRvRR_1q1 _)aha X__XZmah_ _1a )Xu_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a _hXXa_Zh_m_1a aX_ uu)_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRC
M8RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
V`H8RCVm_epB me)h_m
C
oMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RRRRRPOFC#s_00Ns_CCPM
0:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRR#s0N0P_CC2M0RR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"N#0sC0_P0CMRPOFC8sC"
2;RRRRR8CM
RRR
RRRRVRHRe5mpm_Be_ )Bhm) m)_hL2RCMoHRF:RPOD_FsPC_sOFM
CsRRRRRVRHRE5OC_O	FsPCDbNbH2Mo

RRRRRRRORRFsPC_CFPsbDNboHM_N#0sC0_P0CM#R:
RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRRR5H>2R4RR&&#s0N0P_CC2M0RR2
RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5P"FCNsDbMbHo0_#N_s0CMPC0O#RFsPCC28";R
RRCRRMR8
RCRRM
8
CoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
