`ifndef ATCSPI200_CONST_VH
`define ATCSPI200_CONST_VH
`include "ae250_config.vh"
`include "ae250_const.vh"

`define ATCSPI200_PRODUCT_ID		32'h02002046


`ifdef ATCSPI200_AHB_MEM_SUPPORT
	`define ATCSPI200_AHBBUS_EXIST
`elsif ATCSPI200_REG_AHB
	`define ATCSPI200_AHBBUS_EXIST
`endif

`ifdef ATCSPI200_EILM_MEM_SUPPORT
	`define ATCSPI200_EILMBUS_EXIST
`elsif ATCSPI200_REG_EILM
	`define ATCSPI200_EILMBUS_EXIST
`endif

`ifndef ATCSPI200_REG_AHB
	`ifndef ATCSPI200_REG_EILM
		`define ATCSPI200_APBBUS_EXIST
		`ifndef ATCSPI200_REG_APB
			`define ATCSPI200_REG_APB
		`endif
	`endif
`endif

`ifdef ATCSPI200_SPI_ADDR_WIDTH_24
	`define ATCSPI200_SPI_ADDR_WIDTH	24
`else
	`define ATCSPI200_SPI_ADDR_WIDTH	32
`endif
`define ATCSPI200_SPI_ADDR_MSB		(`ATCSPI200_SPI_ADDR_WIDTH - 1)

`ifdef ATCSPI200_ADDR_WIDTH_24
	`define ATCSPI200_HADDR_WIDTH 24
`else
	`define ATCSPI200_HADDR_WIDTH 32
`endif

`define ATCSPI200_HMASTER_BIT 4

`define ATCSPI200_HSPLIT_BIT (1<<`ATCSPI200_HMASTER_BIT)

`ifdef ATCSPI200_AHB_MEM_SUPPORT
	`define ATCSPI200_MEM_SUPPORT
`elsif ATCSPI200_EILM_MEM_SUPPORT
	`define ATCSPI200_MEM_SUPPORT
`endif

`ifdef ATCSPI200_QUADSPI_SUPPORT
	`define ATCSPI200_QUADDUAL_SUPPORT
`elsif ATCSPI200_DUALSPI_SUPPORT
	`define ATCSPI200_QUADDUAL_SUPPORT
`endif

`define ATCSPI200_TXFIFO_WIDTH 32
`define ATCSPI200_RXFIFO_WIDTH 32

`ifdef ATCSPI200_TXFIFO_DEPTH_16W
	`define ATCSPI200_TXFPTR_BITS	5
	`define ATCSPI200_TXFIFO_DEPTH_INF	2'h3
`elsif ATCSPI200_TXFIFO_DEPTH_8W
	`define ATCSPI200_TXFPTR_BITS	4
	`define ATCSPI200_TXFIFO_DEPTH_INF	2'h2
`elsif ATCSPI200_TXFIFO_DEPTH_4W
	`define ATCSPI200_TXFPTR_BITS	3
	`define ATCSPI200_TXFIFO_DEPTH_INF	2'h1
`else
	`define ATCSPI200_TXFPTR_BITS	2
	`define ATCSPI200_TXFIFO_DEPTH_INF	2'h0
`endif

`define ATCSPI200_TXFIFO_DEPTH		(1 << (`ATCSPI200_TXFPTR_BITS - 1))

`ifdef ATCSPI200_RXFIFO_DEPTH_16W
	`define ATCSPI200_RXFPTR_BITS	5
	`define ATCSPI200_RXFIFO_DEPTH_INF	2'h3
`elsif ATCSPI200_RXFIFO_DEPTH_8W
	`define ATCSPI200_RXFPTR_BITS	4
	`define ATCSPI200_RXFIFO_DEPTH_INF	2'h2
`elsif ATCSPI200_RXFIFO_DEPTH_4W
	`define ATCSPI200_RXFPTR_BITS	3
	`define ATCSPI200_RXFIFO_DEPTH_INF	2'h1
`else
	`define ATCSPI200_RXFPTR_BITS	2
	`define ATCSPI200_RXFIFO_DEPTH_INF	2'h0
`endif

`define ATCSPI200_RXFIFO_DEPTH		(1 << (`ATCSPI200_RXFPTR_BITS - 1))

`endif
