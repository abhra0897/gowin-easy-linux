
@ER--=========m==F=FF=========================================FmFF========-
-RR=RB$FbsEHo0BR52jR.4.c-jR4(tHFIMCR1lFHOMO8k0RFsaECOMFFDoB$RFp3,0
83-=-RRRRRRRRRRRRRRRRRRRRRRDqDRosHER0#sCC#s8PC3-
-R====================================================================-=
--
-R_R_RRRRR_R_RRRRR_R_
R--R\\RRRRR/\RRRRRR/RR/RwRrHRDCMCNlR9RRRHbsl$_#ME3P8-
-R\RRRR\R/\R/RR\R/RR/RrRR7OC#s0HbHRFM9WRt4ehR]R7pVOkM0MHFN#DR$EM0C##HRLDHs$Ns
R--R\RRRR\//\RRRR\//RRRRaRrH#lC0bNlR9RRRCakRsqbH.DR6cR4::jjd.jRj
4(-R-RR\RRRRR/R\RRRRR/RRRRRCrPsF#HMRRRRRR9433(n-
-RRRRR/R\RRRRR/R\RRRRRRRRR-
-
R--=========m==F=FF=========================================FmFF========


-------------------------b--NNO	ooCRDNFLD----------------------------
--
ApQ)Yq)RCHCC
;RzR1 HCCC38#0_oDFH4O_43ncN;DDR#
kC RQ 1 3ap7_mBtQ_Qq)aq]3p
p;kR#CQ   371a_tpmQzB_ht1Qh3 7q;pp
q
uBtiq FROlMbFC#M0RRQ1
RRRNs00H0LkC$R#MD_LN_O	L:FGRFLFDMCNRR;
R0RN0LsHkR0C#_$MLODN	F_LGVRFRlBFbCFMMR0#:NRbOo	NC#RHRk0sCR;
R0RN0LsHkR0CLODN	F_LGN_b8H_bM#:R0MsHoR;
R0RN0LsHkR0C#_$MMsFbkRMC:FRLFNDCMR;
R0RN0LsHkR0CGlO_NRb:#H0sM
o;RNRR0H0sLCk0R_GOlRNbFBVRFFlbM0CM#RR:b	NONRoCH"#RD"k0;
RS-N-bOo	NCDRoL#RH
S--#MHoNtDR1R)h:0R#8F_DoRHO:'=R4
';-M-C8DRoL-;
-ObN	CNoR8LF$DRoL-R
-8CMRLoD;-
-----------------------------t-1)-------------------------------------
-
Bumvmhh a1Rt)RR
RuRRmR)a5R
RRRRRRtRR1R)Q:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rt)RR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RM#$_bMFsCkMRRFVtR1):FRBlMbFCRM0H0#Rs;kC
------------------------p--z-a4-----------------------------m
Bvhum Rhap4zaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"";R2
RRRR)uma
R5SRRRR:wRR0FkR8#0_oDFH
O;RRRRRRRRQ:jRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;
0N0skHL0#CR$LM_D	NO_GLFRRFVp4zaRB:RFFlbM0CMRRH#0Csk;0
N0LsHkR0CGlO_NFbRVzRpa:4RRlOFbCFMMH0R#DR"k;0"
-S
-------------------------apz.-R--------------------------
--Bumvmhh azRpa
.RRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"Rj"2R;
RuRRmR)a5R
RRRSRRRRw:kRF00R#8F_Do;HO
RRRSRRRRRQj:MRHR8#0_oDFH
O;RSRRRRRRQ:4RRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRapz.RR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVp.zaRO:RFFlbM0CMRRH#"0Dk"-;
-------------------------apzd----------------------------
--Bumvmhh azRpa
dRRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R""jjR
2;RRRRuam)RR5
RRRSRwRRRF:Rk#0R0D8_FOoH;R
RRRSRRjRQRH:RM0R#8F_Do;HO
RRRSRRRRRQ4:MRHR8#0_oDFH
O;RSRRRRRRQ:.RRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVpdzaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRad:FROlMbFCRM0H"#RD"k0;-
-------------------------pczaR----------------------------B-
mmvuha hRapzcRR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjj";R2
RRRR)uma
R5RSRRRRRRwRR:FRk0#_08DHFoOR;
RRRSRQRRjRR:H#MR0D8_FOoH;R
RRRSRR4RQRH:RM0R#8F_Do;HO
RRRSRRRRRQ.:MRHR8#0_oDFH
O;RSRRRRRRQ:dRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVpczaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRac:FROlMbFCRM0H"#RD"k0;-
-------------------------p6zaR----------------------------B-
mmvuha hRapz6RR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjj";R2
RRRR)uma
R5RSRRRRRRwRR:FRk0#_08DHFoOR;
RRRSRQRRjRR:H#MR0D8_FOoH;R
RRRSRR4RQRH:RM0R#8F_Do;HO
RRRSRRRRRQ.:MRHR8#0_oDFH
O;RSRRRRRRQ:dRRRHM#_08DHFoOR;
RRRSRQRRcRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRa6:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:6RRlOFbCFMMH0R#DR"k;0"
------------------------p--zRan-----------------------------B

mmvuha hRapznRR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjj";R2
RRRR)uma
R5RSRRRRRRwRR:FRk0#_08DHFoOR;
RRRSRQRRjRR:H#MR0D8_FOoH;R
RRRSRR4RQRH:RM0R#8F_Do;HO
RRRSRRRRRQ.:MRHR8#0_oDFH
O;RSRRRRRRQ:dRRRHM#_08DHFoOR;
RRRSRQRRcRR:H#MR0D8_FOoH;R
RRRSRR6RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:nRRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapznRR:ObFlFMMC0#RHRk"D0
";-------------------------z-pa-(R----------------------------
m
Bvhum Rhap(zaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR
2;RRRRuam)RR5
RRRSRwRRRF:Rk#0R0D8_FOoH;R
RRRSRRjRQRH:RM0R#8F_Do;HO
RRRSRRRRRQ4:MRHR8#0_oDFH
O;RSRRRRRRQ:.RRRHM#_08DHFoOR;
RRRSRQRRdRR:H#MR0D8_FOoH;R
RRRSRRcRQRH:RM0R#8F_Do;HO
RRRR6SQRH:RM0R#8F_Do;HO
RRRSRRRRRQn:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRapz(RR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVp(zaRO:RFFlbM0CMRRH#"0Dk"-;
-------------------------apzU-R--------------------------
--
vBmu mhhpaRzRaU
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"2R;
RuRRmR)a5R
RRRSRRRRw:kRF00R#8F_Do;HO
RRRSRRRRRQj:MRHR8#0_oDFH
O;RSRRRRRRQ:4RRRHM#_08DHFoOR;
RRRSRQRR.RR:H#MR0D8_FOoH;R
RRRSRRdRQRH:RM0R#8F_Do;HO
RRRSRRRRRQc:MRHR8#0_oDFH
O;RSRRRRRRQ:6RRRHM#_08DHFoOR;
RRRSRQRRnRR:H#MR0D8_FOoH;R
RRRSRR(RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:URRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapzURR:ObFlFMMC0#RHRk"D0
";-------------------------z-vX-.-----------------------------
m
Bvhum Rhav.zXRR
RRmRu)5aR
RSRRjRQRH:RM0R#8F_Do;HO
RSRR4RQRH:RM0R#8F_Do;HO
RSRRjR1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvX:.RRlBFbCFMMH0R#sR0k
C;-------------------------z-vXp._z-a6-----------------------------B

mmvuha hRXvz.z_pa
6RRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRR1:jRRRHM#_08DHFoOS;
RRRRmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apz6RR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvz.z_pa-n-----------------------------
m
Bvhum Rhav.zX_apznRR
RuRRmR)a5R
SRQRRjRR:H#MR0D8_FOoH;R
SRQRR4RR:H#MR0D8_FOoH;R
SR1RRjRR:H#MR0D8_FOoH;R
SRmRRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.pnzaRB:RFFlbM0CMRRH#0Csk;-
-------------------------v.zX_apz(----------------------------
--
vBmu mhhvaRz_X.p(zaRR
RRmRu)5aR
RSRRjRQRH:RM0R#8F_Do;HO
RSRR4RQRH:RM0R#8F_Do;HO
RSRRjR1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRa(:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.pUza-----------------------------
-
Bumvmhh azRvXp._zRaU
RRRR)uma
R5SRRRRRQj:MRHR8#0_oDFH
O;SRRRRRQ4:MRHR8#0_oDFH
O;SRRRRR1j:MRHR8#0_oDFH
O;SRRRR:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_pa:URRlBFbCFMMH0R#sR0k
C;-------------------------z-vXv._z-XU-----------------------------B

mmvuha hRXvz.z_vX
URRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRR1:jRRRHM#_08DHFoOS;
RRRRmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_XvzURR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvz.z_vX-4n-----------------------------B

mmvuha hRXvz.z_vXR4n
RRRR)uma
R5SRRRRRQj:MRHR8#0_oDFH
O;SRRRRRQ4:MRHR8#0_oDFH
O;SRRRRR1j:MRHR8#0_oDFH
O;SRRRR:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_vXR4n:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.vdzX.----------------------------
--
vBmu mhhvaRz_X.vdzX.RR
RuRRmR)a5R
SRQRRjRR:H#MR0D8_FOoH;R
SRQRR4RR:H#MR0D8_FOoH;R
SR1RRjRR:H#MR0D8_FOoH;R
SRmRRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.vdzX.RR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvzc----------------------------
--
vBmu mhhvaRzRXc
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
SQ:.RRRHM#_08DHFoO
;RSdRQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
S1:4RRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzcRR:BbFlFMMC0#RHRk0sC-;
-------------------------XvzU----------------------------
--
vBmu mhhvaRzRXU
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
SQ:.RRRHM#_08DHFoO
;RSdRQRH:RM0R#8F_Do;HO
QSRcRR:H#MR0D8_FOoH;R
SQ:6RRRHM#_08DHFoOS;
RRQn:MRHR8#0_oDFH
O;S(RQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
S1:4RRRHM#_08DHFoOS;
RR1.:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvX:URRlBFbCFMMH0R#sR0k
C;-------------------------z-vX-4n----------------------------
m
Bvhum Rhav4zXn
RRRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
QSR.RR:H#MR0D8_FOoH;SR
RRQd:MRHR8#0_oDFH
O;ScRQRH:RM0R#8F_Do;HO
QSR6RR:H#MR0D8_FOoH;R
SQ:nRRRHM#_08DHFoOS;
RRQ(:MRHR8#0_oDFH
O;SURQRH:RM0R#8F_Do;HO
QSRgRR:H#MR0D8_FOoH;R
SQR4j:MRHR8#0_oDFH
O;S4RQ4RR:H#MR0D8_FOoH;R
SQR4.:MRHR8#0_oDFH
O;S4RQdRR:H#MR0D8_FOoH;R
SQR4c:MRHR8#0_oDFH
O;S4RQ6RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
RR14:MRHR8#0_oDFH
O;S.R1RH:RM0R#8F_Do;HO
1SRdRR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv4zXnRR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvzd-.--------------------------
--
vBmu mhhvaRz.XdRRR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;S.RQRH:RM0R#8F_Do;HORR
SQ:dRRRHM#_08DHFoOS;
RRQc:MRHR8#0_oDFH
O;S6RQRH:RM0R#8F_Do;HO
QSRnRR:H#MR0D8_FOoH;R
SQ:(RRRHM#_08DHFoOS;
RRQU:MRHR8#0_oDFH
O;SgRQRH:RM0R#8F_Do;HO
QSR4:jRRRHM#_08DHFoOS;
R4Q4RH:RM0R#8F_Do;HO
QSR4:.RRRHM#_08DHFoOS;
RdQ4RH:RM0R#8F_Do;HO
QSR4:cRRRHM#_08DHFoOS;
R6Q4RH:RM0R#8F_Do;HO
QSR4:nRRRHM#_08DHFoOS;
R(Q4RH:RM0R#8F_Do;HO
QSR4:URRRHM#_08DHFoOS;
RgQ4RH:RM0R#8F_Do;HO
QSR.:jRRRHM#_08DHFoOS;
R4Q.RH:RM0R#8F_Do;HO
QSR.:.RRRHM#_08DHFoOS;
RdQ.:HRRM0R#8F_Do;HO
QSR.:cRRRHM#_08DHFoOS;
R6Q.RH:RM0R#8F_Do;HO
QSR.:nRRRHM#_08DHFoOS;
R(Q.RH:RM0R#8F_Do;HO
QSR.:URRRHM#_08DHFoOS;
RgQ.RH:RM0R#8F_Do;HO
QSRd:jRRRHM#_08DHFoOS;
R4QdRH:RM0R#8F_Do;HORR
S1:jRRRHM#_08DHFoOS;
RR14:MRHR8#0_oDFH
O;S.R1RH:RM0R#8F_Do;HO
1SRdRR:H#MR0D8_FOoH;R
S1:cRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzd:.RRlBFbCFMMH0R#sR0k
C;-------------------------p-qz-------------------------------
m
Bvhum RhaqRpz
RRRRht  B)QRR5R
RRRRRRRR7Rq7RR:Q hatR ):j=RRR;
RRRRRRRS1RzA:hRQa  t)=R:R;4R
RRRRRRRR7Rq7A1zRQ:Rhta  :)R=RR.;R
RRRRRRhSR RR:Q hatR ):d=RRR;
RRRRRRRSt: RRaQh )t RR:=c
R;SRRRR RpRQ:Rhta  :)R=;R6
RRRRRRRSzRBuRR:Q hatR ):n=RRR;
RRRRRRRRBR7h:hRQa  t)=R:R;(R
RRRRRRRRzRBuhB7RQ:Rhta  :)R=;RU
RSRRvRRzRpa:hRQa  t)=R:R
g;SRRRRpRqzm_v7: RRaQh )t RR:=jR
RR;R2SR
RRmRu)5aR
1SRz:vRRamzR8#0_oDFH
O;SmRBz:aRRamzR8#0_oDFHSO;
QSRjRR:Q#hR0D8_FOoH;R
SQR4:Q#hR0D8_FOoH;R
SQRd:Q#hR0D8_FOoH;R
SB:QhRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzqpRB:RFFlbM0CMRRH#0Csk;-
--------------------------w-7w-R-----------------------------
m
Bvhum Rha7Rww
RRRRht  B)QRQ5RhRQa:HRL0=R:R''j2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRR:BbFlFMMC0#RHRk0sC-;
-------------------------w-7w- R--------------------------------
m
Bvhum Rha7 wwRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
RRB :hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w RR:BbFlFMMC0#RHRk0sC-;
------------------------71wwR--------------------------------
-
Bumvmhh awR7w
1RRRRRt  h)RQB5hRQQRa:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R1aRR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRw1:FRBlMbFCRM0H0#Rs;kC
----------------------------w7w1- -------------------------------------
m
Bvhum Rha71ww RR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R1aRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw w1RB:RFFlbM0CMRRH#0Csk;-
----------------------w-7w-)R---------------------------------B

mmvuha hRw7w)RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R)1R a:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w)RR:BbFlFMMC0#RHRk0sC-;
-------------------------w-7wR) -------------------------------------B

mmvuha hRw7w)
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
)SR a1 RQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wR) :FRBlMbFCRM0H0#Rs;kC
----------------------------w7wu---------------------------------------
m
Bvhum Rha7uwwRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R u)1: aRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7uwwRB:RFFlbM0CMRRH#0Csk;-
-------------------------7uww -R------------------------------------------
--
vBmu mhh7aRw wuRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R u)1R a:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wu: RRlBFbCFMMH0R#sR0k
C;-----------------------------w7wB-R------------------------------
-
Bumvmhh awR7w
BRRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:BRRlBFbCFMMH0R#sR0k
C;-----------------------------w7wB- R-----------------------------------------
-
Bumvmhh awR7wRB 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw wBRB:RFFlbM0CMRRH#0Csk;-
-------------------------7hwwR----------------------------
--
vBmu mhh7aRwRwh
RRRRht  B)QRQ5RhRQa:HRL0=R:R''j2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:hRRlBFbCFMMH0R#sR0k
C;-----------------w-7wRh ---------------------------------B

mmvuha hRw7wh
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSR RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw whRB:RFFlbM0CMRRH#0Csk;-
----------------------7--w1whR--------------------------------
-
Bumvmhh awR7wRh1
RRRRht  B)QRQ5Rh:QaR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
1SR :aRRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww1RR:BbFlFMMC0#RHRk0sC-;
-------------------------7--w1wh ------------------------------------
--
vBmu mhh7aRw1wh RR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R1aRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw1wh RR:BbFlFMMC0#RHRk0sC-;
----------------------------7hww)--------------------------------
--
vBmu mhh7aRw)whRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R1)  :aRRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww)RR:BbFlFMMC0#RHRk0sC-;
-------------------------w-7w h)R------------------------------------
-
Bumvmhh awR7w h)RR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R1)  :aRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww): RRlBFbCFMMH0R#sR0k
C;----------------------------7hwwu---------------------------------------
m
Bvhum Rha7hwwuRR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S)Ru a1 :hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:uRRlBFbCFMMH0R#sR0k
C;-------------------------w-7w huR--------------------------------------------
-
Bumvmhh awR7w huRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R u)1R a:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whRu :FRBlMbFCRM0H0#Rs;kC
----------------------------w-7wRhB--------------------------------------------
m
Bvhum Rha7hwwBRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:BRRlBFbCFMMH0R#sR0k
C;-----------------------------w7whRB -----------------------------------------
--
vBmu mhh7aRwBwh RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whRB :FRBlMbFCRM0H0#Rs;kC
--------------------------------R7p-----------------------------------------
-
Bumvmhh apR7RR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7RB:RFFlbM0CMRRH#0Csk;-
----------------------7--p- ----------------------------------B

mmvuha hR 7pRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7 RR:BbFlFMMC0#RHRk0sC-;
----------------------------7RpB------------------------------------
m
Bvhum Rha7RpB
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRB7pRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--pRB ------------------------------------
m
Bvhum Rha7 pBRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R Bpq:)RRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7B: RRlBFbCFMMH0R#sR0k
C;-----------------------------u7pR------------------------------------B

mmvuha hRu7pRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RR8#0_oDFH
O;S)Ru a1 RQ:Rh0R#8F_Do;HOSR
StQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:uRRlBFbCFMMH0R#sR0k
C;-----------------------------u7p -R----------------------------------
-
Bumvmhh apR7u
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu7p RR:BbFlFMMC0#RHRk0sC-;
---------------------7--p-hR-----------------------------------------B

mmvuha hRh7pRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7hRR:BbFlFMMC0#RHRk0sC-;
----------------------------7 ph---------------------------------
--
vBmu mhh7aRpRh 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7p RR:BbFlFMMC0#RHRk0sC-;
----------------------------7BphR------------------------------------B

mmvuha hRh7pBRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRhB:FRBlMbFCRM0H0#Rs;kC
----------------------------p-7hRB ------------------------------------
m
Bvhum Rha7Bph RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp hBRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--pRhu------------------------------------
m
Bvhum Rha7uphRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RR8#0_oDFH
O;S)Ru a1 RQ:Rh0R#8F_Do;HOSR
StQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRhu:FRBlMbFCRM0H0#Rs;kC
----------------------------p-7hRu ------------------------------------
m
Bvhum Rha7uph RR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S)Ru a1 RQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7uph RR:BbFlFMMC0#RHRk0sC-;
---------------------zQAw------------------------------------
-
Bumvmhh aARQz
wRRRRRuam)RR5
RSRRR:mRRamzR8#0_oDFH
O;RRRRSRRQ:hRQR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzQAwRR:BbFlFMMC0#RHRk0sC-;
-----------------------------zmAw---------------------------------------
m
Bvhum RhamwAzRR
RRmRu)5aR
RRRRmSRRm:Rz#aR0D8_FOoH;R
RRRRSQRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVRARzw:FRBlMbFCRM0H0#Rs;kC
------------------------------------zaAw---------------------------
m
Bvhum RhaawAzRR
RRmRu)5aR
RRRRRSm:zRma0R#8F_Do;HO
RRRRRSQ:hRQR8#0_oDFH
O;RRRRShm RQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVARaz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFaVRARzw:FRBlMbFCRM0H"#Rm
";
----------------------------AQmz-w------------------------------
-
Bumvmhh amRQARzw
RRRR)uma
R5RRRRSRmR:zRmaRRR#_08DHFoOR;
RSRRQ:mRRmQhz#aR0D8_FOoH;R
RRSRRQ:RRRRQhR#RR0D8_FOoH;R
SRmRR :hRRRQhR#RR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRmwAzRB:RFFlbM0CMRRH#0Csk;-
------------------------------Q--7-7)-------------------------B

mmvuha hR7Q7)RR
RtRR )h Q5BR
jST_QQhaRR:LRH0:'=Rj
';S_T4QahQRL:RH:0R=jR''R
RR;R2SR
RRmRu)5aR
TSRjRR:mRza#_08DHFoOS;
RRT4:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SB:piRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7Q7)RR:BbFlFMMC0#RHRk0sC-;
--------------------------------Q)77B---------------------------
m
Bvhum RhaQ)77BRR
RtRR )h Q5BRRT
Sjh_QQ:aRR0LHRR:=';j'
4ST_QQhaRR:LRH0:'=RjR'
R2RR;RS
RuRRmR)a5R
ST:jRRamzR8#0_oDFH
O;S4RTRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R BpqR):Q#hR0D8_FOoH;SS
RiBp:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ7R)B:FRBlMbFCRM0H0#Rs;kC
-
------------------------------7m7)--------------------
--
vBmu mhhmaR7R7)
RRRRht  B)QR
5RRRRRRRRRapXBim_upRR:LRH0:'=RjR';-j-''H:)#oHMRoC8CkRF00bk;4R''N:wDMDHo8RCoFCRkk0b0RRRRRRRRR
RRRRRRmRBhq1ahQaRhRQa:0R#8F_DoRHO:'=Rj
'RRRRR2
;SRRRRuam)R
5RSRRRRRTj:zRma0R#8F_Do;HOSR
SRTRR4RR:mRza#_08DHFoO
;SSRRRRR7j:hRQR8#0_oDFH
O;SRRRRR74:hRQR8#0_oDFH
O;SRRRRRaX:hRQR8#0_oDFH
O;SRRRRiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR7R7):FRBlMbFCRM0H0#Rs;kC
-
------------------------------7m7)-B---------------------
vBmu mhhmaR7B7)RR
RR RthQ )BRR5
RRRRRRRRBaXpui_m:pRR0LHRR:=';j'R'--j)':HM#Ho8RCoFCRkk0b0';R4w':NHDDMCoR8RoCFbk0kR0RRRRRRRR
RRRRRBRRmah1qRhaQahQR#:R0D8_FOoHRR:='Rj'
RRRRS2;
RRRR)uma
R5SjRTRm:Rz#aR0D8_FOoH;SS
RRT4:zRma0R#8F_Do;HOSR
S7:jRRRQh#_08DHFoOS;
RR74:hRQR8#0_oDFHSO;
aSRXRR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do;HO
BSRp) q:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7R)B:FRBlMbFCRM0H0#Rs;kC
-
--------------------------------------Q--7c 1-----------------------------
--
vBmu mhhQaR7c 1Rt
S )h Q5BR
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)hRR:#H0sM:oR=0R"s"kC
;S2
mSu)5aR
7SSRQ:Rh0R#8F_Do;HO
BSSqApQRQ:Rh0R#8F_Do;HO
)SS a1 RQ:Rh0R#8F_Do;HO
wSSBRpi:hRQR8#0_oDFH
O;SBSup:iRRRQh#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoOS;
SRT.:zRma0R#8F_Do;HO
TSSdRR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71:cRRlBFbCFMMH0R#sR0k
C;
------------------------------------QQe7- m-----------------------------
-
Bumvmhh aeRQQm7 RR
RR RthQ )B
R5S1St)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7RR:Q#hR0D8_FOoH;S
S)  1aRR:Q#hR0D8_FOoH;S
SBQqpARR:Q#hR0D8_FOoH;S
SwiBpRQ:Rh0R#8F_Do;HO
uSSBRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRe Q7mRR:BbFlFMMC0#RHRk0sC-;
---------------------------------7-Q -1U------------------------------------
m
Bvhum RhaQ17 URR
RtRR )h Q5BR
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7 ,)1R a:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;SBSwpui,BRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH;S
ST:(RRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71:URRlBFbCFMMH0R#sR0k
C;
------------------------------------Q--74 1j--------------------------------
--
vBmu mhhQaR74 1jRR
RtRR )h Q5BR
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7 ,)1R a:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;SBSwpui,BRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH;S
ST:(RRamzR8#0_oDFH
O;SUSTRm:Rz#aR0D8_FOoH;S
ST:gRRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71R4j:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------- Q71-4n------------------------------------
vBmu mhhQaR74 1nR
RR RthQ )B
R5RRRRRRRRt 1)hRR:#H0sM:oR=VR"NCD#"R;
RRRRRpRR1h) R#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5R
RRRRRR,R7)  1aRR:Q#hR0D8_FOoH;R
RRRRRRqRBpRQA:hRQR8#0_oDFH
O;RRRRRRRRwiBp,puBiRR:Q#hR0D8_FOoH;R
RRRRRRjRTRm:Rz#aR0D8_FOoH;R
RRRRRR4RTRm:Rz#aR0D8_FOoH;R
RRRRRR.RTRm:Rz#aR0D8_FOoH;R
RRRRRRdRTRm:Rz#aR0D8_FOoH;R
RRRRRRcRTRm:Rz#aR0D8_FOoH;R
RRRRRR6RTRm:Rz#aR0D8_FOoH;R
RRRRRRnRTRm:Rz#aR0D8_FOoH;R
RRRRRR(RTRm:Rz#aR0D8_FOoH;R
RRRRRRURTRm:Rz#aR0D8_FOoH;R
RRRRRRgRTRm:Rz#aR0D8_FOoH;R
RRRRRR4RTjRR:mRza#_08DHFoOR;
RRRRRTRR4:4RRamzR8#0_oDFH
O;RRRRRRRRTR4.:zRma0R#8F_Do;HO
RRRRRRRRdT4Rm:Rz#aR0D8_FOoH;R
RRRRRR4RTcRR:mRza#_08DHFoOR;
RRRRRTRR4:6RRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 4:nRRlBFbCFMMH0R#sR0k
C;
-
----------------------m--1c )-----------------------------
-
Bumvmhh a1Rm R)c
 SthQ )B
R5S1St)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k;C"
RRRRRRRRp]WR#:R0MsHo=R:RN"VD"#C;-R-"k0sCR";"DVN#
C"RRRRRRRRapXBim_upRR:LRH0:'=Rj-'R-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bk
;S2
mSu)5aR
7SSjRR:H#MR0D8_FOoH;S
S7:4RRRHM#_08DHFoOS;
SR7.:MRHR8#0_oDFH
O;SdS7RH:RM0R#8F_Do;HO
aSSX:jRRRHM#_08DHFoOS;
S4aXRH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSwp:iRRRHM#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1):cRRlBFbCFMMH0R#sR0k
C;
--------------------Qme7- m---------------------------------B

mmvuha hRQme7R m
 SthQ )BS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sCS"
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SR7c:MRHR8#0_oDFH
O;S6S7RH:RM0R#8F_Do;HO
7SSnRR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SRST:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVRe Q7mRR:BbFlFMMC0#RHRk0sC-;
-----------------m--1U )---------------------------------
--
vBmu mhhmaR1U )RR
RR RthQ )B
R5RRRRS)t1 :hRRs#0HRMo:"=RV#NDC
";RRRRS)p1 :hRRs#0HRMo:"=R0Csk"R;
RRRRR]RRW:pRRs#0HRMo:"=RV#NDC
";RRRRRRRRapXBim_upRR:LRH0:'=Rj-'R-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bk
RRRR
2;RRRRuam)RR5
RRRRR7RSjRR:H#MR0D8_FOoH;R
RRRRRR4S7RH:RM0R#8F_Do;HO
RRRRRRRSR7.:MRHR8#0_oDFH
O;RRRRRSRR7:dRRRHM#_08DHFoOR;
RRRRR7RScRR:H#MR0D8_FOoH;R
RRRRRSR76:MRHR8#0_oDFH
O;RRRRRSRR7:nRRRHM#_08DHFoOR;
RRRRR7RS(RR:H#MR0D8_FOoH;R
RRRRRRXSajRR:H#MR0D8_FOoH;R
RRaRSX:4RRRHM#_08DHFoOS;
RRRRaRX.:MRHR8#0_oDFH
O;SRRRRdaXRH:RM0R#8F_Do;HO
RSRRBRup:iRRRHM#_08DHFoOS;
RRRR)  1aRR:H#MR0D8_FOoH;R
SRwRRBRpi:MRHR8#0_oDFH
O;RRRRRSRRT:jRRamzR8#0_oDFH
O;RRRRRSRRT:4RRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1):URRlBFbCFMMH0R#sR0k
C;
-------------------- m1)-4j---------------------------------
-
Bumvmhh a1Rm j)4Rt
S )h Q5BR
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)hRR:#H0sM:oR=0R"s"kC
;S2
mSu)5aR
7SSjRR:H#MR0D8_FOoH;S
S7:4RRRHM#_08DHFoOS;
SR7.:MRHR8#0_oDFH
O;SdS7RH:RM0R#8F_Do;HO
7SScRR:H#MR0D8_FOoH;S
S7:6RRRHM#_08DHFoOS;
SR7n:MRHR8#0_oDFH
O;S(S7RH:RM0R#8F_Do;HO
7SSURR:H#MR0D8_FOoH;S
S7:gRRRHM#_08DHFoOS;
SpuBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SwiBpRH:RM0R#8F_Do;HO
TSSRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 4:jRRlBFbCFMMH0R#sR0k
C;
-------------------- m1)-4n---------------------------------B-
mmvuha hR m1)
4nRRRRRht  B)QRR5
RRRRRRRRt 1)hRR:#H0sM:oR=VR"NCD#"R;
RRRRRRRRp 1)hRR:#H0sM:oR=0R"s"kC
RRRR;R2
RRRRmRu)5aR
RRRRRRRRjR7RH:RM0R#8F_Do;HO
RRRRRRRR4R7RH:RM0R#8F_Do;HO
RRRRRRRR.R7RH:RM0R#8F_Do;HO
RRRRRRRRdR7RH:RM0R#8F_Do;HO
RRRRRRRRcR7RH:RM0R#8F_Do;HO
RRRRRRRR6R7RH:RM0R#8F_Do;HO
RRRRRRRRnR7RH:RM0R#8F_Do;HO
RRRRRRRR(R7RH:RM0R#8F_Do;HO
RRRRRRRRUR7RH:RM0R#8F_Do;HO
RRRRRRRRgR7RH:RM0R#8F_Do;HO
RRRRRRRR4R7jRR:H#MR0D8_FOoH;R
RRRRRR7RR4:4RRRHM#_08DHFoOR;
RRRRRRRR7R4.:MRHR8#0_oDFH
O;RRRRRRRRRd74RH:RM0R#8F_Do;HO
RRRRRRRR4R7cRR:H#MR0D8_FOoH;R
RRRRRR7RR4:6RRRHM#_08DHFoOR;
RRRRRRRRuiBpRH:RM0R#8F_Do;HO
RRRRRRRR R)1R a:MRHR8#0_oDFH
O;RRRRRRRRRpwBiRR:H#MR0D8_FOoH;R
RRRRRRRRRRRRRR:TRRamzR8#0_oDFHRO
RRRR2C;
MB8Rmmvuha h;R
RRRRRRRRRR0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 4:nRRlBFbCFMMH0R#sR0k
C;
--------------------7Qm Ypq---------------------------------
--
vBmu mhhQaRmp7 q
YRSht  B)QRR5RBa_1qBaQ_Y7pRH:RMo0CC:sR=2Rj;-R-R4j~.S(
uam)RS5
SR7Q:hRQR8#0_oDFH
O;S7S1aRqu:hRQR8#0_oDFH
O;S S1a:hRRRQh#_08DHFoOS;
Speqz: RRRQh#_08DHFoOS;
SR7m:zRma0R#8F_Do;HO
7SSwRR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7Qm YpqRB:RFFlbM0CMRRH#0Csk;-
------------------ -Qv--------------------------------
--
vBmu mhhQaR 
vRSht  B)Q5S
SW1QhQRZ :0R#soHMRR:="q1vp;p"
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)hRR:#H0sM:oR=0R"s"kC
;S2
mSu)5aR
7SSRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SpvBiH:RM0R#8F_Do;HO
pSSq:tRR0FkR8#0_oDFH
O;S Spq:7RR0FkR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV RQvRR:BbFlFMMC0#RHRk0sC
;
--------------------------------)4qvn-14-------------------------B

mmvuha hRv)q44n1RR
RR RthQ )BRR5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jjRj"2R;
RuRRmR)a5S
S7:mRR0FkR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
SWR) :MRHR8#0_oDFH
O;S7SqRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;SQS7RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n4RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41-.-------------------------
m
Bvhum Rha)4qvnR1.
RRRRht  B)QRQ5Rh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
"RRRRRRRRRRRRR2R;
RuRRmR)a5S
S7:mRR0FkR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
SRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SR7Q:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnR1.:FRBlMbFCRM0H0#Rs;kC
--------------------------------v)q4cn1-------------------------
-
Bumvmhh aqR)v14ncRR
RtRR )h QRB5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RSRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRhRQQ.a_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R;
RRRRRRRRRRRRQahQ_:dRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj
j"RRRRRRRRR2RR;R
RRmRu)5aR
7SSmRR:FRk0#_08DHFoOC_POs0F58dRF0IMF2Rj;SR
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
SRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SR7Q:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnR1c:FRBlMbFCRM0H0#Rs;kC
--------------------------------v)q47n1u-4-------------------------

RRBumvmhh aqR)v14n7Ru4
RRRRht  B)Q5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj";R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S)SW RR:H#MR0D8_FOoH;S
SWRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
S7)qRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;SQS7RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n7Ru4:FRBlMbFCRM0H0#Rs;kC
--------------------------------v)q47n1u-.-------------------------
m
Bvhum Rha)4qvnu17.RR
RtRR )h Q5BRRQQhaR_j:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
SRRRRRQQhaR_4:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj
RRRRRRRRRRRR
2;RRRRuam)RS5
RRRR7:mRR0FkR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
RRRRBRpi:MRHR8#0_oDFH
O;SRRRR W)RH:RM0R#8F_Do;HO
RSRRqRW7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RSRRqR)7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RSRRQR7RH:RM0R#8F_Do_HOP0COF4s5RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRv)q47n1u:.RRlBFbCFMMH0R#sR0k
C;--------------------------------)4qvnu17c------------------------
--
vBmu mhh)aRqnv41c7uRR
RR RthQ )BRR5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RSRRRRRQahQ_:4RR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RRRRRRRRRRRRQRRh_Qa.RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";RRRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R
RRRRRRRRRR;R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH_OPC05FsdFR8IFM0R;j2
BSSp:iRRRHM#_08DHFoOS;
S W)RH:RM0R#8F_Do;HO
WSSq:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S)Rq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SR7Q:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu17cRR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--mnv4-----------------------------B

mmvuha hRv)m4
nRRRRRt  h)RQB5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj";R2
RRRR)uma
R5RRSRRmR7RF:Rk#0R0D8_FOoH;R
SRqRR7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVmR)vR4n:FRBlMbFCRM0H0#Rs;kC



---------------------b--)-mv-------------------------
--Bumvmhh a)Rbm
vRRRRRt  h)RQB5SR
RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SR
SR)RR _q7v m7RL:RH:0R=jR''R;
RRRRR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBSRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRRRRRR
R2RR;R
RRmRu)5aR
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsj.,d2S;
RRRRB,piR,B R mB, R)1R a:MRHR8#0_oDFH
O;SRRRRRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRmb)vRR:BbFlFMMC0#RHRk0sC
;
-----------------------------)-bmgvXR--------------------------------------------B-
mmvuha hRmb)vRXg
RRRRht  B)QR
5RRRRRRRRRA_QaWaQ7]RR:HCM0oRCs:;=g
RRRRRRRRq) 7m_v7: RR0LHR':=j
';RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RRRRRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RR
RR
RRRR
2;RRRRuam)RS5
RRRR7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
RSRRpRBiB,R m,RBR ,)  1aRR:H#MR0D8_FOoH;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFbVR)XmvgRR:BbFlFMMC0#RHRk0sC
;

-

---------------------m-)v----------------------------B

mmvuha hRv)mRR
RR RthQ )BRR5
RSRRQRAaQ_W7Ra]:MRH0CCos=R:4
;SSRRRRq) 7m_v7: RR0LHRR:=';j'
RRRRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRR
RRRRRR2R;
RuRRmR)a5R
SR7RRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SRRRRiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoOR;
RSRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRm:vRRlBFbCFMMH0R#sR0k
C;-----------------------------m-)vRXg---------------------------------------------B

mmvuha hRv)mX
gRRRRRt  h)RQB5RR
RRRRRARRQWa_Q]7aRH:RMo0CC:sR=
g;RRRRRRRR)7 q_7vm RR:LRH0:j=''R;
RRRRRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hRB
RRRRRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRR

R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SpRBiB,R B,m  ,)1, aWR) :MRHR8#0_oDFH
O;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRv)mX:gRRlBFbCFMMH0R#sR0k
C;
-------------------1-u--------------------------------------m
Bvhum Rha1
uRRRRRt  h)RQB5R
SA_QaWaQ7]RR:HCM0oRCs:.=d;-R-RR4,.c,R,,RUR,4nR
d.S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SWa)Q m_v7: RR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SB,piR,B m,B )  1a),W RR:H#MR0D8_FOoH;R
Sq:7RRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRR1u:FRBlMbFCRM0H0#Rs;kC
-
--------------------------u-1X-g--------------------------------------m
Bvhum Rha1guXRR
RR RthQ )BRR5
ASRQWa_Q]7aRH:RMo0CC:sR=
g;S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SWa)Q m_v7: RR0LH_OPC0RFs:j="jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
RiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;R
SB,piR,B m,B )  1a),W RR:H#MR0D8_FOoH;R
Sq:7RRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
RR7Q:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2R

R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRX1ugRR:BbFlFMMC0#RHRk0sC
;

-
---------------------------------1A7u-------------------------------------
--Bumvmhh a7R1u
ARRRRRt  h)RQB5SR
RRRRA_QaWaQ7]R_j:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.R
SRARRQWa_Q]7a_:4RR0HMCsoCR4:=n-;R-,R4RR.,cU,R,nR4,.Rd
RSRR R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
RRRRRRpRAi _1pR_j:HRL0C_POs0FRR:="jjj"R;
RRRRRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"R
RRRRRR2R;
RuRRmR)a5R
SR7RRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SRRRRiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 ARR:H#MR0D8_FOoH;R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRRARRp i1pAq,p i1p:ARRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SR7RRQRR:H#MR0D8_FOoH_OPC05Fsd84RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF1VR7RuA:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------1X7ug-A--------------------------------------m
Bvhum Rha1X7ug
ARRRRRt  h)RQB5SR
RRRRA_QaWaQ7]R_j:MRH0CCos=R:4RU;-g-R,UR4,nRd
RSRRQRAaQ_W7_a]4RR:HCM0oRCs:U=4;-R-RRg,4RU,dSn
RRRR)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSRRRRiAp_p1 _:jRR0LH_OPC0RFs:"=Rj"jj;R
SRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;R
SRBRRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  RaA:MRHR8#0_oDFH
O;SRRRRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRRRRRiAp1q p,iAp1A pRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SRRRRR7Q:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu17XRgA:FRBlMbFCRM0H0#Rs;kC
-
--------------------------u-7A---------------------------------------
m
Bvhum Rha7RuA
RRRRht  B)QRS5
SQRAaQ_W7_a]jRR:HCM0oRCs:n=4;SR
SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;SR
S R)qv7_mj7 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S)RWQ_a v m7jRR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
S)RWQ_a v m74RR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8RC
RSRRRiAp_p1 _:jRR0LH_OPC0RFs:"=Rj"jj;R
RRRRSA_pi1_ p4RR:L_H0P0COF:sR=jR"j;j"
RRRRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
ShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R
RR;R2
RRRR)uma
R5S7SRm7q,m:ARR0FkR8#0_oDFHPO_CFO0s654RI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5j4;n2
RSSBqpi,iBpAB,R Bq, mA,B, qmAB ,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
RSSq,7qqR7A:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;RRRRSpRAip1 qp,Aip1 ARR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RSS7,Qq7RQA:MRHR8#0_oDFHPO_CFO0s654RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRA7uRB:RFFlbM0CMRRH#0Csk;-

-------------------------7--uAXg-------------------------------------
--Bumvmhh auR7XRgA
RRRRht  B)QR
5RSRRRRaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUR
SRARRQWa_Q]7a_:4RR0HMCsoCR4:=U-;R-,RgR
4USRRRRq) 7m_v7R j:HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SR)RR _q7v m74RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSRRRRQW)av _mj7 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
SRWRR) Qa_7vm :4RR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRRRRRA_pi1_ pjRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRRiAp_p1 _:4RR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRR
R2RR;R
RRmRu)5aR
RSRRmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2=R:RMOFP0_#8F_Do_HOP0COFjs5,24U;R
SRBRRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;SRRRRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RSRRQR7qRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;R
RRRRRRpRAip1 qp,Aip1 ARR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RSRRQR7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuAXgRB:RFFlbM0CMRRH#0Csk;



-
---------------------------------1-7u-------------------------------------
-
Bumvmhh a7R1uRR
RtRR )h Q5BRRR
SA_QaWaQ7]R_j:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.R
SA_QaWaQ7]R_4:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.R
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
Rqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds54FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7R1uRR:BbFlFMMC0#RHRk0sC
;
---------------------------------7-1u-Xg-------------------------------------B-
mmvuha hRu17X
gRRRRRt  h)RQB5SR
RaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUd,RnR
SA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4,nRd
)SR _q7v m7RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
RiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
S7:QRRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV1X7ugRR:BbFlFMMC0#RHRk0sCS;

--------------------------------s--1-7u-------------------------------------B-
mmvuha hR7s1uRR
RtRR )h Q5BRRR
SA_QaWaQ7]R_j:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.R
SA_QaWaQ7]R_4:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.R
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A aRH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
S7:QRRRHM#_08DHFoOC_POs0F5Rd48MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVsu17RB:RFFlbM0CMRRH#0Csk;-

---------------------------------7s1u-Xg-------------------------------------B-
mmvuha hR7s1uRXg
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:U=4;-R-RRg,4RU,dSn
RaAQ_7WQa4]_RH:RMo0CC:sR=;4URR--g4,RUd,RnR
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
RRRRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
BSRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  RaA:MRHR8#0_oDFH
O;S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRARRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
7SRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR1X7ugRR:BbFlFMMC0#RHRk0sC
;
---------------------s--)-mv-------------------------
--Bumvmhh a)Rsm
vRRRRRt  h)RQB5SR
RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SR
SR)RR _q7v m7RL:RH:0R=jR''R;
RRRRRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SRBRRpRi,BR ,m,B R1)  :aRRRHM#_08DHFoOR;
RSRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR)Rmv:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------sv)mX-gR--------------------------------------------
vBmu mhhsaR)XmvgRR
RtRR )h Q5BRRR
RRRRRRQRAaQ_W7Ra]:MRH0CCos=R:gR;
RRRRR)RR _q7v m7RL:RH:0R=''j;R
RRRRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
RRRRRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
R
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB,BRm ),R a1 RH:RM0R#8F_Do;HO
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV)RsmgvXRB:RFFlbM0CMRRH#0Csk;

S
-----------------------------7u-------------------------------------
-
Bumvmhh auR7RR
RR RthQ )B
R5SASRQWa_Q]7a_:jRR0HMCsoCR4:=n
;RSASRQWa_Q]7a_:4RR0HMCsoCR4:=n
;RS)SR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)SR _q7v m74RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSWSR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CSWSR) Qa_7vm :4RR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRSpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
ShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R
RR;R2
RRRR)uma
R5S7SRm7q,m:ARR0FkR8#0_oDFHPO_CFO0s654RI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5j4;n2
RSSBqpi,iBpAB,R Bq, mA,B, qmAB ,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
RSSq,7qqR7A:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;RRRRSpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;S7SRQ7q,Q:ARRRHM#_08DHFoOC_POs0F5R468MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7:uRRlBFbCFMMH0R#sR0k
C;
----------------------------X7ug---------------------------------------
vBmu mhh7aRuRXg
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:U=4;-R-RRg,4SU
RaAQ_7WQa4]_RH:RMo0CC:sR=;4URR--g4,RUR
S)7 q_7vm :jRR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
)SR _q7v m74RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)RWQ_a v m7jRR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
RQW)av _m47 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RR
RRRRRR2R;
RuRRmR)a5R
S7,mq7RmA:kRF00R#8F_Do_HOP0COF4s5(FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,24U;R
SBqpi,iBpAB,R Bq, mA,B, qmAB ,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
Rq7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuRXg:FRBlMbFCRM0H0#Rs;kC
-
------------------A--z-wt-------------------------
-
Bumvmhh azRAw
tRRmRu)
a5RRRRS:mRR0FkR8#0_oDFH
O;RRRRS:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVAtzwRB:RFFlbM0CMRRH#0Csk;-
--------------A--z-w1-----------------
--
vBmu mhhAaRzRw1
RRRR)uma
R5RRRRRRRRR:mRR0FkR8#0_oDFH
O;RRRRRRRRR:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVA1zwRB:RFFlbM0CMRRH#0Csk;-
---------------------t-h7----------------
m
Bvhum RhatRh7
RRRR)uma
R5RRRRSRRt:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVhRt7RR:BbFlFMMC0#RHRk0sC-;
--------------------e-BB---------------------
--
vBmu mhheaRB
BRRRRRuam)RR5
RSRRR:eRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRBeBRB:RFFlbM0CMRRH#0Csk;

S-----------------1-mB-w--------------------------
-
Bumvmhh a1RmB
wRRRRRt  h)RQB5R
RRRRRR)Rw 7T_Q:eRR0HMCsoCRR:=gRnR-~-.gFn,MRD$CMPCRlMk
RRRR
2;RRRRuam)RS5
RRRRmm1Bz:aRR0FkR8#0_oDFH
O;RRRRRRRRmm1Bzjadvm:Rz1aRap7_mBtQ;R
RRRRRR1RmBR h:hRQR71a_tpmQRB
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRBm1wRR:BbFlFMMC0#RHRk0sC
;
-----------------eQh---------------------------------B

mmvuha hReQhRR
RRmRu)5aR
RRRRmSRRm:Rz#aR0D8_FOoH;R
RRRRSQRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRh:eRRlBFbCFMMH0R#sR0k
C;
-

-----------------Bm1Z----------------------------B

mmvuha hRBm1ZRR
RtRR )h Q5BR
RRRRRRRR w)TQ_7eRR:HCM0oRCs:4=RjRjR-~-.4,.UF$MDRCCPMkRMlR
RR;R2
RRRR)uma
R5SRRRRBm1mSza:kRF00R#8F_Do;HO
mSS1hB SQ:RhaR17m_ptSQBRR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVmZ1BRB:RFFlbM0CMRRH#0Csk;


-----------------eap7Q1_A-zw--------------------------------
m
Bvhum Rhaa7pe1A_QzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH;R
RRRRRRARQRQ:Rh0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFReap7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1A_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------eap7m1_A-zw--------------------------------
m
Bvhum Rhaa7pe1A_mzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRm:ARRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpRae_71mwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFReap7m1_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------p-ae_71awAz---------------------------------B

mmvuha hReap7a1_A
zwRRRRuam)RR5
RSRRRRmR:zRmaRRR#_08DHFoOR;
RSRRRRmA:zRma0R#8F_Do;HO
RRRRRRSQ:RRRRQhR#RR0D8_FOoH;R
SRRRRmR h:hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFaVRp1e7_zaAwRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpRae_71awAzRB:RFFlbM0CMRRH#"Rm,m;A"
-
--------------a--p1e7_AQmz-w------------------------------
--
vBmu mhhaaRp1e7_AQmzRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSQRmA:hRQmRza#_08DHFoOR;
RRRRRRRRQ:mRRmQhz#aR0D8_FOoH;R
RRSRRRRQR:hRQRRRR#_08DHFoOS;
RRRRRhm RQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVa7pe1m_QARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1m_QARzw:FRBlMbFCRM0H"#RQRm,Q"mA;-

---------------- 7pe1A_Qz-w------------------------------
--
vBmu mhh aRp1e7_zQAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFHRO
RRRRR2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFV 7pe1A_Qz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMF VRp1e7_zQAwRR:BbFlFMMC0#RHR,"QR"QA;-

---------------- 7pe1A_mz-w------------------------------
--
vBmu mhh aRp1e7_zmAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRmRRARR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7m1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_mz:wRRlBFbCFMMH0R#mR",ARm"
;
-----------------e p7a1_A-zw--------------------------------
m
Bvhum Rha 7pe1A_azRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSm:ARRamzR8#0_oDFH
O;RRRRRQSRRRR:QRhRR0R#8F_Do;HO
RSRRmRR :hRRRQhR#RR0D8_FOoH
RRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpR e_71awAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRe p7a1_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------p- e_71QzmAw--------------------------------
-
Bumvmhh apR e_71QzmAwR
RRmRu)5aR
RRRRmSRRRR:mRzaR0R#8F_Do;HO
RRRRQSRm:ARRmQhz#aR0D8_FOoH;R
RRRRRRQRRmRR:Qzhma0R#8F_Do;HO
RRRRRRSQ:RRRRQhR#RR0D8_FOoH;R
SRRRRmR h:hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGF VRp1e7_AQmz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMF VRp1e7_AQmz:wRRlBFbCFMMH0R#QR"mQ,Rm;A"



------------------------vQQu_zQAw------------------------------------m
Bvhum RhavQQu_zQAwR
RRmRu)5aR
RRRRRRRR]Rm,pRm,ARmRm:Rz#aR0D8_FOoH;R
RRRRRRQRRmQ,Rm:ARRmQhz#aR0D8_FOoH;R
RRRRRRQRR,ARQRQ:Rh0R#8F_Do;HO
RRRRRRRR Rmhm,R ,hAR)]1 :hRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFvVRQ_uQQwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRuvQQA_Qz:wRRlBFbCFMMH0R#QR"mQ,Rm;A"
-
R---------------------v--Q_uQQwAz_-]1---------------------------------
--Bumvmhh aQRvuQQ_A_zw]R1
RRRRuam)RR5
RRRRRRm]:zRma0R#8F_Do;HO
RRRRQRRRQ:Rh0R#8F_Do;HO
RRRRQRRARR:Q#hR0D8_FOoH
RRRR;R2
MRC8mRBvhum ;ha
RRRR0RN0LsHkR0C#_$MLODN	F_LGVRFRuvQQA_Qz]w_1RR:BbFlFMMC0#RHRk0sCR;
RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFvVRQ_uQQwAz_R]1:FRBlMbFCRM0H"#RQQ,RA
";
-R---------------------vQQu_zQAwu_p-------------------------------------B
Rmmvuha hRuvQQA_Qzpw_uR
RRuRRmR)a5R
RRRRRRRRRm:pRRamzR8#0_oDFH
O;SRRSRRmA:zRma0R#8F_Do;HOSR
RRRRRRRRRQRR:Q#hR0D8_FOoH;R
SSQRRARR:Q#hR0D8_FOoH
RRRR;R2
MRC8mRBvhum ;ha
RRRR0RN0LsHkR0C#_$MLODN	F_LGVRFRuvQQA_Qzpw_uRR:BbFlFMMC0#RHRk0sCR;
RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFvVRQ_uQQwAz_Rpu:FRBlMbFCRM0H"#RQQ,RA
";
-R----------------------Q-vumQ_A-zw-------------------------------------R-
Bumvmhh aQRvumQ_A
zwRRRRR)uma
R5RRRRRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRRmRRARR:mRza#_08DHFoOR;
RRRRRRRRR:QRRRQh#_08DHFoOS;
RRSRQ:ARRRQh#_08DHFoOR;
RRRRRRRRR7vm p1 RQ:Rh0R#8F_Do
HORRRRR
2;R8CMRvBmu mhh
a;RRRRR0N0skHL0#CR$LM_D	NO_GLFRRFVvQQu_zmAwRR:BbFlFMMC0#RHRk0sCR;
RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFvVRQ_uQmwAzRB:RFFlbM0CMRRH#"Rm,m;A"
-
--------------------------d-QBm_QA-zw-----------------------------
--
vBmu mhhQaRdQB_mwAzRR
RRmRu)5aR
RRRRRSmRm:RzRaRR8#0_oDFH
O;RRRRSRQm:hRQmRza#_08DHFoOR;
RRRRSRQR:hRQRRRR#_08DHFoOS;
RRRRv m71R p:hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ_dBQzmAwRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVdRQBm_QARzw:FRBlMbFCRM0H"#RQ;m"
S

R-
--------------------------q-u7U74-------------------------------------
--Bumvmhh aqRu7U74
oSSCsMCH
O5SRSRR)Rq :tRR0LHRR:=';j'-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SRRRRAt) RL:RH:0R=jR''
;RSRSRRmR1)R t:HRL0=R:R''j;S
SRRRRq_771RzA:HRL0=R:R''j;R
RRRRRRRRRRqRu7)7_ a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-Rh1YB1,qY
hBRRRRRRRRRRRRAp1 _7vm RR:LRH0:'=R4-'R-4R""#:RE0HV,jR""b:RNDsNDRCDHkMb03RA
RSRR;R2
RRRRRRR
RRRRRRRRsbF0S5
SRRRR:qRRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SRRRR:ARRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SRRRR q1pRR:H#MR0D8_FOoH;S
SRRRRBB ,p)i, a1 RH:RM0R#8F_Do;HO
RSSR1RRQA,1QRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SRRRR11m,A:mRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0FjR2
RSRR2 ;
hB7Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqRu7U74RB:RFFlbM0CMRRH#0Csk;-

-------------------------u--qg77-------------------------------------
--Bumvmhh aqRu7
7gRRRRRRRRoCCMs5HO
RSSRqRR)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SRRRR A)tRR:LRH0:'=RjR';
RSSR1RRmt) RL:RH:0R=jR''S;
SRRRR7q7_A1zRL:RH:0R=jR''R;
RRRRRRRRRuRRq_77)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-YR1hqB,1BYh
RRRRRRRRRRRR A1pm_v7: RR0LHRR:='R4'-"-R4R":#VEH0",RjR":bNNsDDDCRbHMkA0R3R
SR2RR;R
RRRRRRRR
RSRRb0FsRS5
SRRRR:qRRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
SRRRRARR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
RSSRqRR1R p:MRHR8#0_oDFH
O;SRSRR RB,iBp,1)  :aRRRHM#_08DHFoOS;
SRRRR,1Q1RAQ:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SRRRR,1m1RAm:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;SRSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0sR5U8MFI0jFR2R
SR2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7uq7:gRRlBFbCFMMH0R#sR0k
C;
----------------------------pvzaggX-------------------------------------m
Bvhum Rhavazpg
XgSCSoMHCsOS5
SRRRR q)tRR:R0LHRR:=';j'RR--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CSRSRR)RA :tRRHRL0=R:R''j;S
SRRRRm_za)R t:LRRH:0R=jR''S;
SRRRRuuQ  _)tRR:R0LHRR:=';j'
RSSRqRR1hQt_t) RR:RLRH0:'=Rj
';SRSRR1RAQ_th)R t:LRRH:0R=jR''R;
RRRRRRRRR1RRm)q_ :tRRHRL0=R:R''j;SR
SRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
RRRR2
;
RRRRSsbF0
R5SRSRR,Rq1RQq:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SRRRR1A,Q:ARRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
SRRRRqt1QhA,R1hQtRH:RM0R#8F_Do;HO
RRRRRRRRRRRR q1p1,A :pRRRHM#_08DHFoOS;
SRRRRRB :MRHR8#0_oDFH
O;SRSRRpRBiRR:H#MR0D8_FOoH;S
SRRRR)  1aRR:H#MR0D8_FOoH;S
SRRRR7amzRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj;R
RRRRRRRRRRmR1qm,1ARR:FRk0#_08DHFoOC_POs0F58URF0IMF2Rj
RSRR;R2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpgRXg:FRBlMbFCRM0H0#Rs;kC
-
--------------------------z-vpUa4X-4U-------------------------------------
-
Bumvmhh azRvpUa4X
4URRRRoCCMs5HO
qSS)R t:LRRH:0R=jR''-;R-'RRjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SAt) RR:RLRH0:'=Rj
';SzSma _)tRR:R0LHRR:=';j'
uSSQ_u )R t:LRRH:0R=jR''S;
SQq1t)h_ :tRRHRL0=R:R''j;S
SAt1Qh _)tRR:R0LHRR:=';j'
RRRRRRRRq1m_t) RR:RLRH0:'=Rj
';SzSvp)a_ a1 _7vm RR:#H0sM:oR=1R"Y"hBRR--1BYh,1RqY
hBS
2;
FSbs50R
qSS,q1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
ASS,A1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
qSS1hQt,1RAQRth:MRHR8#0_oDFH
O;RRRRRRRRqp1 , A1pRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
7SSmRza:kRF00R#8F_Do_HOP0COFds56FR8IFM0R;j2
RRRRRRRRq1m,A1mRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazp44UXURR:BbFlFMMC0#RHRk0sC
;
----------------------------vazpddnXn---------------------------------------
vBmu mhhvaRzdpannXd
CSoMHCsOS5
S q)tRR:R0LHRR:=';j'RR--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CS)SA :tRRHRL0=R:R''j;S
Smjza_t) RR:RLRH0:'=Rj
';SzSma)4_ :tRRHRL0=R:R''j;S
Su Qu_t) RR:RLRH0:'=Rj
';S1SqQ_th)R t:LRRH:0R=jR''S;
SQA1t)h_ :tRRHRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
S:qRRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
S:ARRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
SQq1tRh,At1QhRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
7SSmRza:kRF00R#8F_Do_HOP0COF(s54FR8IFM0R
j2S
2; Rh7Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzdpannXdRB:RFFlbM0CMRRH#0Csk;-

-------------------------v--zqpapnzdX-4U-------------------------------------B-
mmvuha hRpvzazqpd4nXUo
SCsMCH
O5S)Sq :tRRHRL0=R:R''j;-R-RjR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
ASS)R t:LRRH:0R=jR''S;
S B)tRR:R0LHRR:=';j'
mSSz)a_ :tRRHRL0=R:R''j;S
Su Qu_t) RR:RLRH0:'=Rj
';S1SqQ_th)R t:LRRH:0R=jR''S;
SQA1t)h_ :tRRHRL0=R:R''j;R
RRRRRRBRqBqpm7 _)t:jRR0LHRR:=';j'
RRRRRRRRBqBp7mq_t) 4RR:LRH0:'=Rj
';RRRRRRRR1_mq)R t:HRL0=R:R''j;R
RRRRRRzRvppaqzXdn4vU_mR7 :MRH0CCos=R:R-j;-dj:nUG4R-+/RRB;4B:qBR/j+nRdG;4URR.:d4nGURR+BQq1
RRRRRRRRqB_717_z:ARR0LHRR:=';j'-'-RjR':N;88R4R''#:RkSL
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2R;
R
RRSsbF0
R5SRSq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSA:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;SRSB:MRHR8#0_oDFHPO_CFO0sd56RI8FMR0Fj
2;S1SqQ,thRQA1tRh,qpBBmRq7:MRHR8#0_oDFH
O;S SBRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
S1BqQRR:H#MR0D8_FOoH_OPC05Fs68cRF0IMF2Rj;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;S
SBmq1RF:Rk#0R0D8_FOoH_OPC05Fs68cRF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpqdpznUX4RB:RFFlbM0CMRRH#0Csk;R
RR-R
-------------------------v--zqpa7p7qzX4U4-U--------------------------------------m
Bvhum Rhavazpqq77pUz4X
4USMoCCOsH5S
Sq j)tRR:LRH0:'=Rj-';-jR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
ASSjt) RL:RH:0R=jR''
;RS4Sq)R t:HRL0=R:R''j;S
SA 4)tRR:LRH0:'=Rj
';S)SB :tRR0LHRR:=';j'
mSSz)a_ :tRR0LHRR:=';j'
uSSQju _t) RL:RH:0R=jR''S;
SuuQ )4_ :tRR0LHRR:=';j'
qSS1hQtj _)tRR:LRH0:'=Rj
';S1SAQjth_t) RL:RH:0R=jR''S;
SQq1t_h4)R t:HRL0=R:R''j;S
SAt1Qh)4_ :tRR0LHRR:=';j'
qSSBmBpq)7_ Rtj:HRL0=R:R''j;S
SqpBBm_q7)4 tRL:RH:0R=jR''R;
RRRRR1RRm)q_ :tRR0LHRR:=';j'
ASS_7q7_A1zRL:RH:0R=jR''R;R-'-RjR':N;88R''4:kR#LS
SB7_q7z_1ARR:LRH0:'=Rj
';SzSvp7aq7zqp44UXUm_v7: RR0HMCsoCRR:=j-;-jU:4GR4U+R/-44UGU/R+-;RBR:R4RBqB/+jRRG4U4+UR/4-RUUG4;:R.44UGU/R+-UR4GR4U+qRB1SQ
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5SjSq,Rq4:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SjSA,RA4:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SQS1qQ,1ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SBRR:H#MR0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R
RRRRRR1RqQ,thAt1QhRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RRRRRRRR q1p1,A :pRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRRqRB1:QRRRHM#_08DHFoOC_POs0F5R6c8MFI0jFR2R;
RRRRRqRRBmBpq:7RRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R
RRRRRRmR1qm,1ARR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
S1BqmRR:FRk0#_08DHFoOC_POs0F5R6c8MFI0jFR22
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvza7q7q4pzUUX4RB:RFFlbM0CMRRH#0Csk;-

-------------------------v--zqpapUz4X-4U-------------------------------------B-
mmvuha hRpvzazqp44UXUo
SCsMCH
O5S)Sq :tRR0LHRR:=';j'-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SAt) RL:RH:0R=jR''
;RS)SB :tRR0LHRR:=';j'
7SS)R t:HRL0=R:R''j;R
RRRRRRzRma _)tRR:LRH0:'=Rj
';SQSuu) _ :tRR0LHRR:=';j'
qSS1hQt_t) RL:RH:0R=jR''S;
SQA1t)h_ :tRR0LHRR:=';j'
7SS1hQt_t) RL:RH:0R=jR''S;
SBqBp7mq_t) jRR:LRH0:'=Rj
';SBSqBqpm7 _)t:4RR0LHRR:=';j'
ASS_7q7_A1zRL:RH:0R=jR''R;R-'-RjR':N;88R''4:kR#LS
SB7_q7z_1ARR:LRH0:'=Rj
';SzSvppaqzX4U4vU_mR7 :MRH0CCos=R:R-j;-qj:BjB/R-+/RG4U4+UR/B-R;:R4q/BBj/R+-UR4GR4U+qRB1RQ;.4:RUUG4R-+/R+7RR1BqQS;
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5SRSq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSA:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;S,SBR:7RRRHM#_08DHFoOC_POs0F5R6d8MFI0jFR2R;
RRRRRqRR1hQt,1RAQRth:MRHR8#0_oDFH
O;RRRRRRRRBQq1RH:RM0R#8F_Do_HOP0COF6s5cFR8IFM0R;j2
RRRRRRRRBqBp7mq,Q71t:hRRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;S
SBmq1RF:Rk#0R0D8_FOoH_OPC05Fs68cRF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpq4pzUUX4RB:RFFlbM0CMRRH#0Csk;-

-------------------------q--pcz67------------------------------------
--Bumvmhh apRqz76c
CSoMHCsOS5
RRRRqt) RL:RH:0R=jR''-;R-''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CRRRRRRRRAt) RL:RH:0R=jR''S;
RRRRqt1Qh _)tRR:LRH0:'=Rj
';SRRRRQA1t)h_ :tRR0LHRR:=';j'
RSRRBRqBqpm7 _)tRR:LRH0:'=Rj
';SRRRRamz_t) RL:RH:0R=jR''S;
RRRRA7_q7z_1ARR:LRH0:'=Rj-';-''j:8N8;4R''k:#LR
SRBRR_7q7_A1zRL:RH:0R=jR''R;
RRRRRqRRp_z7v m7RH:RMo0CC:sR=;Rj-:-jq/BBj/R+-RRA+R/-q4;R:BqB/+jR/A-RRB+Rq;1QRq.:R-+/R+ARR1BqQS;
Szqp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-h1YBq,R1BYh
RRRR
2;RRRRb0FsRS5
RRRRqRR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRARR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRB: RRRHM#_08DHFoOS;
RRRRBRpi:MRHR8#0_oDFH
O;SRRRR1)  :aRRRHM#_08DHFoOS;
RRRRqt1Qh1,AQRth:MRHR8#0_oDFH
O;SRRRRBqBp7mqRH:RM0R#8F_Do;HO
RSRRqRB1:QRRRHM#_08DHFoOC_POs0FRc56RI8FMR0Fj
2;SRRRRz7maRR:FRk0#_08DHFoOC_POs0FRd56RI8FMR0Fj
2;SRRRR1BqmRR:FRk0#_08DHFoOC_POs0FRc56RI8FMR0FjR2
R2RR;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzqp6Rc7:FRBlMbFCRM0H0#Rs;kC
-
------------------------------p-up------------------------
--Bumvmhh apRupR
RR RthQ )BR5
RRRRRRRRRRRRwiBpQ:hRR)1aQRht:"=R43jjjR";-s-VCCJkMRO$F0VREOCRDM	H5
v2RRRRRRRRRRRRRe7 QRB :aR1)tQhRR:="4tWh"-.;-R-"4tWh"-4,W"t4.h-"t,"W-4hc"",thW4-,n"RW"t4gh-"t,"W)4h-,c""4tWhg)-"t,"W-4h.,A""4tWhA-c"t,"W)4h-"cA,W"t4nh- ,1""4tWh -g1"",thW4) -g1"",thW41"-.,W"t4-h1.
B"RRRRRRRRRRRRRh7Y_QQ7e _1pRR:1Qa)h:tR=VR"NCD#"-;-0Csk:1Q7 Rp;V#NDC7:QQ1e_ Rp
RRRRRRRRRRRRQe7Q_p1 RH:RMo0CC:sR=;Rj-M-QbRk08HHP8RCsQe7Q,:Rj4:,4.333nnd:cR3R4c~n
RRRRRRRRRRRRYR7hA_w7_Qe1R p:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRARw7_Qe1R p:MRH0CCos=R:R-j;-CwC8OLN	HR8PCH8sARw7,QeR:Rj4:,4.333nnd:c43R~
ncRRRRRRRRRRRRRh7Y_Qm7e _1pRR:1Qa)h:tR=VR"NCD#"-;-0Csk:1m7 Rp;V#NDC7:mQ1e_ Rp
RRRRRRRRRRRRme7Q_p1 RH:RMo0CC:sR=;RU-/-.c//U4dn/.U/c//ncUgj/n4/4../4UR
RRRRRRRRRRuRR1_7q1R p:aR1)tQhRR:="jjjj-";-R
RRRRRRRRRR7RRY7h_qh_ R1:Rah)Qt=R:RN"VD"#C;0--s:kCuq17RRFs7Yza7FqRs7RwqV;RNCD#:qR7_p1 
RRRRRRRRRRRRzR7aqY7_p1 R1:Rah)Qt=R:Rj"4j;j"-R-
RRRRRRRRRRRRBmpizwa_aQ_7)RR:LRH0:'=R4R';-B-RpzimaHRVM0CRkMMHoHR8s0COH3FMR''4RDFM$RR
RRRRRRRRRRRRBmpiz_auw7a_Q:)RR0LHRR:=';4'RR--'R4'F$MD
RRRRRRRRRRRRpRBiamz_Y7p_ 1auRR:HCM0oRCs:j=R;-R-R4j,,c.,
RRRRRRRRRRRRpRBiamzup_7Ya_1 :uRR0HMCsoCRR:=j-;R-,Rj4
,.
RRRRRRRRRRRRpRBiamz71d_):BRR)1aQRht:"=RBmpiz;a"-C-#D0CORP8HdkRF00bk,pRBiamzusRFRiBpm
zaRRRRRRRRRRRRRiBpw1A_ :pRR)1aQRht:"=RHCM0sDMN"R;
RRRRRRRRRRRRBmpizAa_Y1uq1RR:1Qa)h:tR=VR"NCD#"R;
RRRRRRRRRRRRBmpiz_auAqYu1:1RR)1aQRht:"=RV#NDC
";RRRRRRRRRRRRRiBpm7za_uAYqR11:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRpRBiamz7)_1BRR:1Qa)h:tR=BR"pzima-";-D#CCRO08RHPFbk0kR0,RiBpmuzaRRFsBmpizRa
RRRRRRRRRRRR7_Yh1e7Q_p1 RH:RMo0CC:sR=RR.-.-R~U4.,DFM$PRCCMMRkRl
RRRRRRRRRRRR
RSRRRRR2R;
RuRRm5)a
RRRRRRRRRRRRpRBiRQh:hRQR8#0_oDFH
O;RRRRRRRRRRRRRiBpw:ARRRQh#_08DHFoO':=j
';RRRRRRRRRRRRR1Q7 :pRRRQM#_08DHFoOC_POs0F586RF0IMF2Rj;R
RRRRRRRRRRwRRA 71pRR:Q#MR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
RRRRRRRRRRRR7Rm1R p:MRQR8#0_oDFHPO_CFO0sR568MFI0jFR2R;
RRRRRRRRRRRR)  1aRR:H#MR0D8_FOoH:j=''R;
RRRRRRRRRRRR)  1aR_u:MRHR8#0_oDFH=O:';j'
RRRRRRRRRRRR R)1_ aQHR:M0R#8F_Do:HO=''j;R
RRRRRRRRRR)RR a1 _:1RRRHM#_08DHFoO=R:';j'
RRRRRRRRRRRR1Ru7wq,7RpY:MRQR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;
RRRRRRRRRRRR7Yza7:qRRRQM#_08DHFoOC_POs0F58dRF0IMF2Rj;R
RRRRRRRRRRpRRmRBi:zRma0R#8F_Do;HO
RRRRRRRRRRRRpRBiamzRm:Rz#aR0D8_FOoH;R
RRRRRRRRRRBRRpzima:7RR0FkR8#0_oDFH
O;RRRRRRRRRRRRRiBpmuzaRF:Rk#0R0D8_FOoH;R
RRRRRRRRRRBRRpzimaR7d:kRF00R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRupRR:BbFlFMMC0#RHRk0sC
;
-----------------p7p---------------------------------m
Bvhum Rha7
ppRRRRt  h)5QB
RRRRRRRRp7p_)wmB: RR0HMCsoCRR:=j-;-4V:RFCsORODF	MRN8FRO8RC;jO:RF/8CD	FORMoCC0sNCV8RsRFl7RppDbFF
RRRRRRRRe7Q_p1 RL:RH:0R=4R''-;-jF,MsDlNRODF	FRl8RC;4N,V#D0RFRO	lCF8
RSRRmRB7B 1q:pRR)1aQRht:"=Rj"jj;j--jj4R4jjR444Rj4jRj44R44jR4R4
RRRRR1RRB_qp :hRR)1aQRht:"=R0Csk"0--s,kCV#NDCR
RR;R2
RRRR)umaR5
RRRRRBRRphiQ:RQh#_08DHFoO':=j
';RRRRRRRR1uam:MRQR8#0_oDFH=O:';j'
RRRRRRRR1)  :aRRRQM#_08DHFoO':=j
';RRRRRRRRzhu7BphaRQ:RM0R#8F_Do:HO=''j;R
RRRRRRmRpB:iRRamzR8#0_oDFH
O;RRRRRRRR1ua Rm:Rz#aR0D8_FOoH_OPC05Fs(FR8IFM0R
j2RRRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:pRRlBFbCFMMH0R#sR0k
C;
--------------------------------iBp7-Qe-------------------------m
Bvhum RhaB7piQRe
RtRR )h Q
B5SRRRRQR7em_v7: RR)1aQRht:"=R.R";-"-R.R","6d3"",RcR",",6"R""U5""U,DmM$kR#bsbF0RC8HoMRI-4Mng	/	S2
RRRRR)t1 :hRR)1aQRht:"=RV#NDC-"R-VR"NCD#"",R0Csk"R
SR2RR;R
RRmRu)
a5RRRRRRRRRp]BiRQh:hRQR8#0_oDFH
O;SRRRR R)1h aRQ:Rh0R#8F_Do;HO
RSRRBRRqApQRQ:RM0R#8F_Do;HO
RSRRBRRpzimaRR:mRza#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVB7piQ:eRRlBFbCFMMH0R#sR0k
C;S-
------------------------------]-7B- h------------------------------------
vBmu mhh7aR]hB 
RRRR)uma
R5SpRBiamzRm:Rz#aR0D8_FOoH;SS
RRB :hRQR8#0_oDFHSO;
BSRphiQRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VR]hB RB:RFFlbM0CMRRH#0Csk;
R
-----------------------------p-7pY7p-------------------------------------
--Bumvmhh apR7pY7p
RRRRht  B)Q5R
RRRRRRpR7ph_Q1R p:HRL0=R:R''j;-R-':j'LN$b#l#RF,8CR''4:#RkCDR8DC_8DRN$ODCD
RRRRRRRRY7p_t1QhRR:LRH0:'=RjR';-'-Rj'':+R',R''4:-R''R
RRRRRRpR7Y7_qKRR:HCM0oRCs:j=RRj--~6.6,DR8$H_#ojM=RD:8$8_N[8;RD#$_H=oM4-:R.+6n8_D$NR8[
RRRR
2;RRRRuam)5R
RRRRRRpR7p 1auRR:Q#hR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRRRRRRiBpQQh:h0R#8F_Do;HO
RRRRRRRR)7Q,qpm7vh,m:e RRQM#_08DHFoOR;
RRRRRBRRpzimaRR:mRza#_08DHFoOR;
RRRRRwRRpRqt:zRma0R#8F_Do
HORRRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRppp7YRR:BbFlFMMC0#RHRk0sC
;R



-----------------------------p-wq.1]6-ni-------------------------------------B-
mmvuha hRqwp16].nRi
RuRRm5)a
RRRRRRRR7Xq)RR:Q#hR0D8_FOoH_OPC05FsnFR8IFM0R;j2
RRRRRRRR7Yq)RR:Q#hR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
RRRRRRRR,X Y1 , h:QR8#0_oDFH
O;RRRRRRRR7RQh:hRQR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2;RRRRRRRR 1)q ),umht,e)1a:hRQR8#0_oDFH
O;RRRRRRRR7amzRm:Rz#aR0D8_FOoH_OPC05Fsd84RF0IMF2Rj
RRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVw1pq]n.6iRR:BbFlFMMC0#RHRk0sCR;RR
R



R
--------------------------------B-71------------------------------------B-
mmvuha hR17B
RRRRht  B)QRS5
S17B_7vm RR:#H0sM:oR=)R"Qh1QtR"RRB--p,ijB4pi,iBp.p,Bitd,he7,B)B,Qh1Qtq,wphpQtp,Bitj_hB7,p_ije,BBB4pi_7th,iBp4B_eBp,Bit._hB7,p_i.e,BBBdpi_7th,iBpdB_eB2
S;u
SmR)a5S
SBjpiRQ:Rh0R#8F_Do;HO
BSSpRi4:hRQR8#0_oDFH
O;SpSBi:.RRRQh#_08DHFoOS;
SiBpdRR:Q#hR0D8_FOoH;S
SB1pi :pRRRQh#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S1w pm )BRQ:Rh0R#8F_Do;HO
BSSpzimaRR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR17BRB:RFFlbM0CMRRH#0Csk;RRRR-

-----------------------------7--T-B ------------------------------------
vBmu mhh7aRT
B RRRRuam)RS5
RiBpmRza:zRma0R#8F_Do;HOSR
SB: RRRQh#_08DHFoO
;SSpRBiRQh:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVTR7B: RRlBFbCFMMH0R#sR0kRC;R
RRR
RR
-
--------------------------p-wq41].-Ui-----------------------------m
Bvhum Rhaw1pq]U4.iR
RRmRu)
a5RRRRRRRRq)77RQ:Rh0R#8F_Do_HOP0COF4s5cFR8IFM0R;j2
RRRRRRRRh7QRQ:Rh0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRR,B1qm , RR:Q#hR0D8_FOoH;R
RRRRRRBRup:iRRRQh#_08DHFoOR;
RRRRRuRR),mt1q ),1vq QR:h0R#8F_Do;HO
RRRRRRRR)Qw )h, a1 he,h1:a)RRQh#_08DHFoOR;
RRRRR7RRmRza:zRma0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRRQaAaRR:mRza#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVw1pq]U4.iRR:BbFlFMMC0#RHRk0sCR;RR
R
-----------------------------B-vz---------------------------------------
vBmu mhhvaRBRz
RuRRm5)a
RRRRRRRRpwBiRR:Q#hR0D8_FOoH;R
RRRRRRmRu)  1a:hRRRQh#_08DHFoOR;
RRRRR1RRY 1)1h aRQ:Rh0R#8F_Do;HO
RRRRRRRRB)a1B)Bp:iRRRQh#_08DHFoOR;
RRRRRQRRmu XmuzazRam:zRma0R#8F_Do_HOP0COF4s56FR8IFM0R;j2
RRRRRRRR QmXzumaauz Rhm:zRma0R#8F_Do_HOP0COF4s56FR8IFM0R;j2
RRRRRRRR QmXhuQuQzaRQ:Rh0R#8F_Do_HOP0COF4s56FR8IFM0R;j2
RRRRRRRR)zqaXja7:mRRamzR8#0_oDFH
O;RRRRRRRRzaq)47aXmRR:mRza#_08DHFoOR;
RRRRRzRRqj)aA7qzaiQBRm:Rz#aR0D8_FOoH;R
RRRRRRqRz)Aa4qaz7QRBi:zRma0R#8F_Do;HO
RRRRRRRR)zqaXj)7:QRRRQh#_08DHFoOR;
RRRRRzRRq4)a)QX7RQ:Rh0R#8F_Do;HO
RRRRRRRRaQhvQmhaRm):zRma0R#8F_Do;HO
RRRRRRRRXva]1)  Rah:zRma0R#8F_Do;HO
RRRRRRRRq1)v7jq7:)RRamzR8#0_oDFHPO_CFO0s.54RI8FMR0Fj
2;RRRRRRRR1v)qj W)hRR:mRza#_08DHFoOC_POs0F58dRF0IMF2Rj;R
RRRRRR)R1qWvj7qqaRm:Rz#aR0D8_FOoH_OPC05Fsd84RF0IMF2Rj;R
RRRRRR)R1qBvj1RR:mRza#_08DHFoOR;
RRRRR1RR)jqv)a7qqRR:H#MR0D8_FOoH_OPC05Fsd84RF0IMF2Rj;R

RRRRRaRRqw)tp]q1j ]1pRR:mRza#_08DHFoOR;
RRRRRaRRqw)tp]q1j7]q7:)RRamzR8#0_oDFHPO_CFO0sU5.RI8FMR0Fj
2;RRRRRRRRatq)w1pq]aj])1qhRm:Rz#aR0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RRRRRRRR)aqtqwp1]]jWa)Q RR:mRza#_08DHFoOR;
RRRRRaRRqw)tp]q1jQ]1Z: RRamzR8#0_oDFHPO_CFO0sR5.8MFI0jFR2R;
RRRRRaRRqw)tp]q1jz]A)R1a:zRma0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;RRRRRRRRatq)w1pq]uj])Rma:zRma0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRatq)w1pq] jvvaqa)RR:mRza#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRRqRa)ptwqj1]  X)TRR:mRza#_08DHFoOR;
RRRRRaRRqw)tp]q1jq]v1)a Rm:Rz#aR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRR)aqtqwp1]]jWa7qqRR:mRza#_08DHFoOC_POs0F5Rd48MFI0jFR2R;
RRRRRaRRqw)tp]q1jq]v1mapB:iRRamzR8#0_oDFH
O;RRRRRRRRatq)w1pq])j] Yq7vRzX:zRma0R#8F_Do;HO
RRRRRRRR)aqtqwp1]]jq z1)RR:mRza#_08DHFoOR;
RRRRRaRRqw)tp]q1jz]W1R ):zRma0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRatq)w1pq])j]7qqaRQ:Rh0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRR)aqtqwp1]]j) z1)RR:Q#hR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RRRRRRRR)aqtqwp1]]j)u 1RQ:Rh0R#8F_Do;HO
RRRRRRRR)aqtqwp1 ]jX1) uRR:Q#hR0D8_FOoH;R
RRRRRRqRa)ptwqj1]]q) 7zYmaRR:Q#hR0D8_FOoH;R

RRRRRaRRq )tX]uj1R p:zRma0R#8F_Do;HO
RRRRRRRR)aqtu Xj7]q7:)RRamzR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2;RRRRRRRRatq) jXu]qa)h:1RRamzR8#0_oDFHPO_CFO0sR548MFI0jFR2R;
RRRRRaRRq )tX]ujWa)Q RR:mRza#_08DHFoOR;
RRRRRaRRq )tX]uj1 QZRm:Rz#aR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RRRRRRRR)aqtu Xjz]A)R1a:zRma0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;RRRRRRRRatq) jXu]mu)aRR:mRza#_08DHFoOC_POs0F58dRF0IMF2Rj;R
RRRRRRqRa)Xt u jvvaqa)RR:mRza#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRRqRa)Xt uXj )R T:zRma0R#8F_Do;HO
RRRRRRRR)aqtu Xjq]v1)a Rm:Rz#aR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRR)aqtu Xj7]WqRaq:zRma0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRR)aqtu Xjq]v1mapB:iRRamzR8#0_oDFH
O;RRRRRRRRatq) jXu]q) 7zYvXRR:mRza#_08DHFoOR;
RRRRRaRRq )tX]ujq z1)RR:mRza#_08DHFoOR;
RRRRRaRRq )tX]ujW z1)RR:mRza#_08DHFoOC_POs0F58dRF0IMF2Rj;R
RRRRRRqRa)Xt u)j]7qqaRQ:Rh0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRR)aqtu Xj ])qm7Yz:aRRRQh#_08DHFoOR;
RRRRRaRRq )tX]uj)u 1RQ:Rh0R#8F_Do;HO
RRRRRRRR)aqtu Xj) X R1u:hRQR8#0_oDFH
O;RRRRRRRRatq) jXu]1)z :)RRRQh#_08DHFoOC_POs0F58.RF0IMF2Rj;R

RRRRRQRRh QaX]uj)a7qqRR:mRza#_08DHFoOC_POs0F5Rd48MFI0jFR2R;
RRRRRQRRh QaX]uj)7 qYRR:mRza#_08DHFoOR;
RRRRRQRRh QaX]uj)u 1Rm:Rz#aR0D8_FOoH;R
RRRRRRhRQQXa uXj )u 1Rm:Rz#aR0D8_FOoH;R
RRRRRRhRQQXa u)j]z)1 Rm:Rz#aR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RRRRRRRRQQhau Xj ]1pRR:Q#hR0D8_FOoH;R
RRRRRRhRQQXa uqj]7R7):hRQR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2;RRRRRRRRQahQ jXu]qa)h:1RRRQh#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRRhRQQXa uWj]) QaRQ:Rh0R#8F_Do;HO
RRRRRRRRQQhau XjQ]1Z: RRRQh#_08DHFoOC_POs0F58.RF0IMF2Rj;R
RRRRRRhRQQXa uAj]za)1RQ:Rh0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;RRRRRRRRQahQ jXu]mu)aRR:Q#hR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRQQhau Xjvv q)aaRQ:Rh0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;RRRRRRRRQahQ jXu  X)TRR:Q#hR0D8_FOoH;R
RRRRRRhRQQXa uvj]q 1a)RR:Q#hR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRQQhau Xj7]WqRaq:hRQR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2;RRRRRRRRQahQ jXu]1vqaBpmiRR:Q#hR0D8_FOoH;R
RRRRRRhRQQXa uqj]z)1 RQ:Rh0R#8F_Do;HO
RRRRRRRRQQhau Xjz]W1R ):hRQR8#0_oDFHPO_CFO0sR5d8MFI0jFR2
;
RRRRRRRRqauAq )tXuu.1Aa)Rm:Rz#aR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRAquatq) .Xuumu)aRR:mRza#_08DHFoOC_POs0F58.RF0IMF2Rj;R
RRRRRRuRqA)aqtu X. u1pRR:mRza#_08DHFoOR;
RRRRRqRRuqAa)Xt u .uhpqA RR:mRza#_08DHFoOR;
RRRRRqRRuqAa)Xt uq.u7R7):zRma0R#8F_Do_HOP0COF4s54FR8IFM0R;j2
RRRRRRRRAquatq) .XuuQW)a: RRamzR8#0_oDFH
O;RRRRRRRRqauAq )tXuu.Wa7qqRR:mRza#_08DHFoOC_POs0F5Rd48MFI0jFR2R;
RRRRRqRRuqAa)Xt u).u7qqaRQ:Rh0R#8F_Do_HOP0COFds54FR8IFM0R;j2
RRRRRRRRAquatq) .Xuuq) 7:YRRRQh#_08DHFoOR;
RRRRRqRRuqAa)Xt u1.up)e )RR:Q#hR0D8_FOoH;R

RRRRRvRRa X)vRqu:hRQR8#0_oDFHPO_CFO0sR5d8MFI0jFR2
;
RRRRRRRR71quWR7m:zRma0R#8F_Do;HO
RRRRRRRRu7q1mW7 :hRRamzR8#0_oDFH
O;RRRRRRRR7aqu7:mRRamzR8#0_oDFH
O;RRRRRRRR7Kquahqt1:WRRamzR8#0_oDFH
O;RRRRRRRR7hqua 7mhRR:mRza#_08DHFoOR;
RRRRR7RRqWu17vQa1RR:Q#hR0D8_FOoH;R
RRRRRRqR7uQa7RQ:Rh0R#8F_Do;HO
RRRRRRRRu7qh1a)aRR:Q#hR0D8_FOoH;R
RRRRRRqR7uB1WpBiaiRR:Q#hR0D8_FOoH;R

RRRRRaRRuaQz) qB7qqaRm:Rz#aR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRQauzqa)BW 1mRR:mRza#_08DHFoOR;
RRRRRaRRuaQz) qBBRpi:zRma0R#8F_Do;HO
RRRRRRRRqwp1)] )RR:Q#hR0D8_FOoH;R
RRRRRRpRwqQ1]h:aRRRQh#_08DHFoOR
RR2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzvBRB:RFFlbM0CMRRH#0Csk;RRRR-

-----------------------------Az1.uj_]-Y--------------------------------------m
Bvhum Rhaz.1Aj]_uYR
RR RthQ )BR5
RRRRRRRRRRRR7qqaA4z1nR_U:HRL0=R:R''j;-R-1CCDOR0#LIC0CRCMUMRN8nR4R0LHR08NNsR0NVM#C
s#RRRRRRRRRRRRRuq7_Au) :hRR0LHRR:=';j'R --MDNLC8#/HL#NDRC#0RECqR7uuLsFCFROlsbNNs0F
RRRRRRRRRRRR Ra1va_mR7 :HRL0C_POs0FRR:=Xj"jj"jj;k--#RC8VRFs00C#HRMoNRM88kCLoMoHokRbs#bFCR
RRRRRRRRRR]RR1e7)4RR:LRH0:'=RjR';-H-]o#ERb8CCRH8sPNCR8#[k0MlC0u3RD#CNCFROMOMC0FR0RVjRFMsRFNslDbRFC0sNH
FMRRRRRRRRRRRRR7]1)Rej:HRL0=R:R''j;R
RRRRRRRRRRBRRp1i_ :pRR0LHRR:=';j'-D-BFRO	#sFkO#CRCODC0MHFRo#HM3NDR0jRFCR#D0COR0CGCNsMDDROFRO	bPsFH88CRRL$0RECO#s$0RNDOMFMCCO08MRFRhXQ,mRXzRa34FR0RD#CCRO0HCM0sDMNRFODOb	RsHFP8RC8FQMRhpaBiFRbsR0
RRRRRRRRRRRRvRR:L_H0P0COF:sR="RXjjjj"-;-vHR8PCH8sMRHbRk08NN0R0LH#R
RRRRRRRRRRhRRRL:RHP0_CFO0s=R:R4X"jj4jj-";-8hRH8PHCHsRM0bkR08NNHRL0R#
RRRRRRRRRRRRBRR:L_H0P0COF:sR="RXjjjj"-;-B0FMsRFDOsENobCRkRlbOsksCRM0HkMb0NR80LNRH,0#RRH0#bkbF#s0RFVsljRdk5qRjRj20nFRjRkq5244
RRRRRRRRRRRRmRwBm_pB:iRR0LHRR:='-j'-Rj:pimBRRH#oCCMsCN08$RLRpupRODF	CR800COFRs34p:RmRBiHN#RD$IN#HREoNE5D$IN#FRDO
	2
RRRRRSRRRRR2R;
RuRRm5)a
RRRRRRRRa7qqamzRm:Rz#aR0D8_FOoH_OPC05Fs486RF0IMF2Rj;R
RRRRRRXRa)7 qYRR:mRza#_08DHFoOR;
RRRRR)RRXaqBQRe :zRma0R#8F_Do;HO
RRRRRRRRe)Xp:7RRamzR8#0_oDFH
O;RRRRRRRR)pXe7:]RRamzR8#0_oDFH
O;RRRRRRRRBRpi:zRma0R#8F_Do;HO
RRRRRRRR )X)))mRm:Rz#aR0D8_FOoH;R
RRRRRRQRpha 1qRa :zRma0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;RRRRRRRR7:uRRmQhz#aR0D8_FOoH;R
RRRRRRvR7RQ:RhamzR8#0_oDFH
O;RRRRRRRR7qqaQ:hRRRQh#_08DHFoOC_POs0F5R468MFI0jFR2R;
RRRRRaRRX7epRQ:Rh0R#8F_Do;HO
RRRRRRRReaXpR7]:hRQR8#0_oDFH
O;RRRRRRRR)  1aRR:Q#hR0D8_FOoH;R
RRRRRRzR11hu 7:vRRRQh#_08DHFoOR;
RRRRRXRRB1e) :pRRRQh#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRR Ra) v1pRR:Q#hR0D8_FOoH;R
RRRRRRuRmv m7RQ:Rh0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;
RRRRRRRR1]ma17QRm:Rz#aR0D8_FOoH;R
RRRRRR7RQ7RQt:zRma0R#8F_Do;HO
RRRRRRRRuq7uR)A:zRma0R#8F_Do;HO
RRRRRRRRuq71Rh1:zRma0R#8F_Do;HO
RRRRRRRR11 17epRm:Rz#aR0D8_FOoH;R
RRRRRRARezp1e7RR:mRza#_08DHFoOR;
RRRRR)RRXR7u:zRma0R#8F_Do;HO
RRRRRRRR7)XvRR:mRza#_08DHFoOR;
RRRRR)RRXe)BRm:Rz#aR0D8_FOoH;R
RRRRRR7RQupzpz:uRRRQh#_08DHFoOR;
RRRRR7RRuRu7:hRQR8#0_oDFH
O;RRRRRRRR77vuRQ:Rh0R#8F_Do;HO
RRRRRRRRqB])Atez:1RRRQh#_08DHFoOR;
RRRRR7RRQ]1Bqe)tARz1:hRQR8#0_oDFH
O;RRRRRRRRaQXAaz1awhw RQ:Rh0R#8F_Do;HO
RRRRRRRRAaXQaa1z wwh:]RRRQh#_08DHFoOR;
RRRRRaRRXh hRQ:Rh0R#8F_Do;HO
RRRRRRRR7aXq:aRRRQh#_08DHFoOR;
RRRRRaRRXj1 RQ:Rh0R#8F_Do;HO
RRRRRRRRpw11)1 QRqp:hRQR8#0_oDFH
O;RRRRRRRRp Ai):)RRamzR8#0_oDFH
O;RRRRRRRRB)pi7:YRRamzR8#0_oDFH
O;RRRRRRRRQBhap:iRRRQh#_08DHFoOR;
RRRRRQRR7RR:Qzhma0R#8F_Do;HO
RRRRRRRRzeA1RR:Qzhma0R#8F_Do;HO
RRRRRRRRX) aRR:Qzhma0R#8F_Do;HO
RRRRRRRRhXQRQ:Rh0R#8F_Do;HO
RRRRRRRRzXmaRR:Qzhma0R#8F_Do;HO
RRRRRRRRiBpcuUjq:7RRamzR8#0_oDFH
O;RRRRRRRRaa 1RQ:Rh0R#8F_Do;HO
RRRRRRRRq1Bhamz4RR:mRza#_08DHFoOR;
RRRRR1RRBmqhzRa.:zRma0R#8F_Do;HO
RRRRRRRRq1BhamzdRR:mRza#_08DHFoOR;
RRRRR1RRBmqhzRac:zRma0R#8F_Do;HO
RRRRRRRRq1Bhamz6RR:mRza#_08DHFoOR;
RRRRR1RRBmqhzRan:zRma0R#8F_Do;HO
RRRRRRRRq1BhiBpRQ:Rh0R#8F_Do;HO
RRRRRRRRq1BhR h:hRQR8#0_oDFH
O;RRRRRRRR1hBqv m7RQ:Rh0R#8F_Do;HO
RRRRRRRR a)1h aRQ:Rh0R#8F_Do;HO
RRRRRRRRq1Bh4QhRQ:Rh0R#8F_Do;HO
RRRRRRRRq1Bh.QhRQ:Rh0R#8F_Do;HO
RRRRRRRRq1BhdQhRQ:Rh0R#8F_Do;HO
RRRRRRRRq1BhcQhRQ:Rh0R#8F_Do;HO
RRRRRRRRq1Bh6QhRQ:Rh0R#8F_Do;HO
RRRRRRRRq1BhnQhRQ:Rh0R#8F_Do
HO
RRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVz.1Aj]_uYRR:BbFlFMMC0#RHRk0sCR;RRRR
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRV1RzA_.juR]Y:FRBlMbFCRM0H"#R7Ru,7Rv,QR7,e1Az, R)XRa,Xamz,QRXh
";RRRR
----------------------------q--7-B--------------------------------------m
Bvhum Rhaq
7BSht  B)Q5S
Sew) _R h:HRL0=R:R''j;-R-jH,8#DNLCR->N_8OPVCs=BeBX4;R,MRCNCLD-F>OMoVHk8sCRRL$bNNslCC0s)Re 1w_ Sp
S e)w _1pRR:L_H0P0COF:sR="RXj"jj-j-jjB,eBRX;j,j4dcc/je5*B2BX;4Rjj4,d/5cj*BeBXR2;j,44.cg/je5*B2BX;jR4j(,./5cj*BeBXR2;4,j4.c./je5*B2BX;4R4jj,./5cj*BeBXR2;4,44VlsFRRQmuRq7ew) 
2SS;R
RRmRu)
a5RRRRRRRRB:]RRRQh#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRRRRR R1pRR:Q#hR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
RRRRRRRRiBp,,u71RmB:hRQR8#0_oDFH
O;RRRRRRRRew) RQ:Rh0R#8F_Do;HO
RRRRRRRRB mRm:Rz#aR0D8_FOoH;R
RRRRRR7RqmRza:zRma0R#8F_Do_HOP0COF4s54FR8IFM0R
j2RRRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFqVR7:BRRlBFbCFMMH0R#sR0k
C;S0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVqR7B:FRBlMbFCRM0H"#RBR],ew) "S;

M
C8FROlMbFC#M0;RRRR







