-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRR:1RR08NMNRs8ep]7RM1$0#ECHu#RNNO	o
C#-R-RRRRRRRRRR:RRRhR5z)v QAB_Qza_ht1QhR 7b	NONRoC8DCON0sNH2FM
R--RRRRRRRRRRRR:-
-RpRRHNLssR$RRR:Ra#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRRR:R#L$lFODHN$DDRlMNCQ8R 3  
R--RRRRRRRRRRRR:-
-R7RRCDPCFsbC#R:RqCOODsDCN]Re7ap-BN,RMQ8R R  u(4jnFRWsM	HosRtF
kb-R-RRRRRRRRRR:RR
R--RkRus#bFCRRR:aRRERH#b	NONRoC8HCVMRC#MCklsRHO0C$b#MRN8sRNHl0ECO0HRMVkOF0HM-#
-RRRRRRRRRRRRRR:RsVFRCk#R0IHE$R#MC0E#RH#0DFF#e3RNCDk#VRFRb0$CQRAa _eB)am
R--RRRRRRRRRRRR:NRRsHCRMs0Cb0sCCN8R#MRk#MHoCM8RkClLsH#RMCRPOs0FRsVFl-3
-RRRRRRRRRRRRRR:RCaERVDC0#lF0HRL0#RHRC0sN80CRRN#0RECl0F#Ro#HMHHVO0NMR0LH3-
-RRRRRRRRRRRRRR:Ra#EHRObN	CNoRMOF0MNH#PRFCFsDN88CRHNs0CEl0RHOFsbCNs0F#MRF
R--RRRRRRRRRRRR:0RREACRQea_ mBa)$R0bRC3aRECb	NONRoCNFD#RMOF0MNH#-
-RRRRRRRRRRRRRR:RkV#Ck0DR$RbCOPFMCHs#FRM#VOkM0MHF#O,RD	FOR08CCHO0F-M
-RRRRRRRRRRRRRR:RMVkOF0HMR#,NRM8FC0Es0RkH0DH$kRVMHO0F3M#
R--RRRRRRRRRRRR:-
-RRRRRRRRRRRRRR:RQNVRMN$RslokCRM00NFRRMVkOF0HM#RHRMNRkRDDNNss$N,RRDMkDsRNs
N$-R-RRRRRRRRRR:RRR#RHR0sCkCsM8CR5GbOC0MHF#H,RVMRN$N,RsMCRF80CR8HMH8PHkDND$
23---
-RRRhCF0RRRRRRR:RHaE#NRbOo	NCNRl$CRLR8lFHCVH8FR0ROHMDCk8R8N8HF0HMRND8NN0
R--RRRRRRRRRRRR:sRRCHJksRC8L0$RF#FD,kRL00RHR#lk0MRHRRMFIRN$OMENo0CRE-C
-RRRRRRRRRRRRRR:R0CGCNsMDMRH0VCsN#OCRRFs#kHlDHN0FLMRCPENHRFsF0VRE-C
-RRRRRRRRRRRRRR:R#8CObsH0MHF30RQRRH#blCsHH##LRDC0NFR8O8RFCllMR0#N/M8F-s
-RRRRRRRRRRRRRR:R0N0skHL0RC#00FREbCRNNO	o8CRCNODsHN0F,M#R0LkR0MFRR0FOMENo-C
-RRRRRRRRRRRRRR:RRFs8CCD0NCRMF$RsHHoMRNDDCHM#VRFRC0ERObN	CNoRO8CDNNs0MHF3-
-RRRRRRRRRRRRRR:RaRECb	NONRoCL$F8R$lNRRLCOMENoRC8F$MDRRHMNFOOsM8NOICRH
0E-R-RRRRRRRRRR:RRRER0CCR0sRl#FBVRD#NkCnR4RRFV0#EHRN#0Ms8N8-3
-RRRRRRRRRRRR
R:---R-----------------------------------------------------------------
---f-R)HCP#MHF:.R4.fjR
R--f07NC.:Rj-jUj4c-j(R4::4nj+gRjjgdRE5ak4,RjbRqsjR.jRU2f-
-R--------------------------------------------------------------------b

NNO	ohCRz)v QAB_Qza_ht1QhR 7HR#
RMOF#M0N0FRBbH$)ohE0FO0HCRR:1Qa)h:tR=R
RRBR"Fsb$H0oERj.jU RQ R 3qRDDsEHo0s#RCs#CP3C8"
;
R-R-R:Q8Rdq3
VRRk0MOHRFM"R+"5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFvs5qvXQzpv5'hp t,a]Rp)' aht]42-RI8FMR0Fj
23R-R-R#)Ck:D0R8q8#IR0FhRz1hQt P7RCFO0s0#RERN0lRN$LFCRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8q:R3
d)RkRVMHO0F"MR+p"5RA:RQea_ mBa));RRA:RQRa2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFps5'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Rl1HHsDNRR0FqR3dIsECCRR)HN#RRCFMR0LHR0LH_OPC0
Fs
-RR-8RQ:3RqdRp
RMVkOF0HM+R""R5p:QRAa);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1HHlDRNs0qFR3IdRECCsRHpR#RRNFRMCLRH0zQh1t7h 
R
R-Q-R8q:R3R6
RMVkOF0HM+R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFps5'hp t-a]4FR8IFM0R3j2
-RR-CR)#0kD:8Rq8N#RMhRz1hQt P7RCFO0sp,R,HRI0NERRMMF-oMCNP0HChRQa  t)),R3R

RR--QR8:q
3nRkRVMHO0F"MR+5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR0LH_OPC05Fs) 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k0q:R8R8#NFRMMC-MoHN0PQCRhta  R),pI,RHR0ENzMRht1QhR 7P0COFRs,)
3
R-R-============================================================================
R
R-Q-R8q:R3Rg
RMVkOF0HM-R""pR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:hRz1hQt v75qvXQzpv5'hp t,a]Rp)' aht]42-RI8FMR0Fj
23R-R-R#)Ck:D0RL1k0OsN00#RIzFRht1QhR 7P0COFRs#00ENR$lNRRLCF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:q)3g
VRRk0MOHRFM"5-"pRR:A_Qaea BmR);)RR:A2QaR0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR0LH_OPC05Fsp 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR1lNHDsFR0Rgq3RCIEs)CRRRH#NMRFCHRL0hRz1hQt 
7
R-R-R:Q8Rgq3pR
RVOkM0MHFR""-5:pRRaAQ;RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RHDlHN0sRF3RqgERICRsCp#RHRFNRMLCRHz0Rht1Qh
 7
-RR-8RQ:3Rq4R4
RMVkOF0HM-R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFps5'hp t-a]4FR8IFM0R3j2
-RR-CR)#0kD:kR1LN0sOR0#NFRMMC-MoHN0PQCRhta  R),)V,RsRFlNzMRht1QhR 7P0COFRs,p
3
R-R-R:Q8R4q3.R
RVOkM0MHFR""-RR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s'5)pt ha4]-RI8FMR0Fj
23R-R-R#)Ck:D0RL1k0OsN0N#RMhRz1hQt P7RCFO0s),R,sRVFNlRRMMF-oMCNP0HChRQa  t)p,R3R

R=--=========================================================================
==
-RR-8RQ:3Rq4R6
RMVkOF0HM*R""pR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5'5ppt ha)]+'hp t-a]482RF0IMF2Rj3R
R-)-RCD#k0u:RCFsVsRl#0RECl0kDHHbDOHN0FFMRbNCs0MHFRRFM0RIFzQh1t7h ROPC0#Fs
-RR-RRRRRRRRER0Nl0RNb$RFH##LRD$LFCRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8q:R3
4(RkRVMHO0F"MR*5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR0LH_OPC05Fs5pp' aht]'+ppt ha4]-2FR8IFM0R3j2
-RR-CR)#0kD:kRvDb0HD#HCRRNMzQh1t7h ROPC0,FsRRp,IEH0RMNRFMM-C0oNH
PCR-R-RRRRRRRRRaQh )t ,3R)RH)R#FROMsPC0RC80NFRMhRz1hQt P7RCFO0sVRF
-RR-RRRRRRRRQR1Zp R'hp tRa]LFCVslCRkHD0bODHNF0HM
3
R-R-R:Q8R4q3UR
RVOkM0MHFR""*RR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s)55'hp t+a]) 'ph]ta-R428MFI0jFR2R3
RR--)kC#DR0:v0kDHHbDCN#RMhRz1hQt P7RCFO0s),R,HRI0NERRMMF-oMCNP0HCR
R-R-RRRRRRQRRhta  R),pp3RRRH#OPFMCCs08FR0RRNMzQh1t7h ROPC0RFsFRV
RR--RRRRRRRR1 QZRp)' aht]CRLVCFsRDlk0DHbH0ONH3FM
R
R-=-==========================================================================R=
R
--R-R-Rahm Q:RVCR#O8FMRoNskMlC0#RHRsxCFFRVs/R""bRFC0sNFRs,NCR#PHCs0D$RCDPC
-RR-RRRRRRRF VR)))mRRH#Hk##C
83
-RR-8RQ:3Rq.R4
RMVkOF0HM/R""pR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5pp' aht]R-48MFI0jFR2R
R-)-RCD#k07:RH8PHCN#RMhRz1hQt P7RCFO0sp,R,$RLRFNM0sECR1zhQ th7CRPOs0F,3R)
R
R-Q-R8q:R3
.dRkRVMHO0F"MR/5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR0LH_OPC05Fsp 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#MRNR1zhQ th7CRPOs0F,,RpRRL$NFRMMC-MoHN0PQCRhta  R),)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:qc3.
VRRk0MOHRFM"R/"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5p)' aht]R-48MFI0jFR2R
R-)-RCD#k07:RH8PHCN#RRMMF-oMCNP0HChRQa  t)p,R,$RLRRNMzQh1t7h ROPC0,FsR
)3R-R-RRRRRRRRRRQVhmm_wQ_Aap152RR>) 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rp)' aht]
3
R-R-============================================================================
-RR-R
R-h-Rm:a RRQV#FCOMN8RslokCRM0Hx#RCRsFVRFs"lsC"bRFC0sNFRs,NCR#PHCs0D$RCDPC
-RR-RRRRRRRF VR)))mRRH#Hk##C
83
-RR-8RQ:3Rq.R(
RMVkOF0HMsR"CRl"5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COF)s5'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"RlsCRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0s
#3
-RR-8RQ:3Rq.Rg
RMVkOF0HMsR"CRl"5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsNRM8)#RHRRN
RR--RRRRRRRRM-FMMNCo0CHPRaQh )t 3R
R-R-RRRRRRQRRVmRh__mwA1Qa5R)2>'Rppt haR],skC#DH0R#sR0kNMO0RC80pFR'hp t3a]
R
R-Q-R8q:R3
djRkRVMHO0F"MRs"ClRR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRH)R#MRNR1zhQ th7CRPOs0FR8NMRHpR#
RNR-R-RRRRRRRRRMMF-oMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0F) 'ph]ta3R

R=--=========================================================================
==R-R-
-RR-mRhaR :Q#VRCMOF8sRNoCklMH0R#CRxsVFRF"sRl"F8RCFbsFN0sN,RRP#CC0sH$CRDP
CDR-R-RRRRRFRRV)R )Rm)HH#R#C#k8
3
R-R-R:Q8Rdq3dR
RVOkM0MHFRF"l85"Rp),RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"plRF8)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#
3
R-R-R:Q8Rdq36R
RVOkM0MHFRF"l85"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR0LH_OPC05Fsp 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpFRl8"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRM)8R
-RR-RRRRRRRR#RHRMNRFMM-C0oNHRPCQ hat3 )
-RR-RRRRRRRRVRQR_hmmAw_Q5a1)>2RRpp' aht]s,RCD#k0#RHRk0sM0ONC08RF'Rppt ha
]3
-RR-8RQ:3RqdRn
RMVkOF0HMlR"FR8"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:HRL0C_POs0F5p)' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsC)#RHRRNMzQh1t7h ROPC0RFsNRM8pR
R-R-RRRRRRHRR#RRNM-FMMNCo0CHPRaQh )t 3R
R-R-RRRRRRQRRVmRh__mwA1Qa5Rp2>'R)pt haR],skC#DH0R#sR0kNMO0RC80)FR'hp t3a]
R
R-=-==========================================================================R=
RR--QR8:qg3d
VRRk0MOHRFMV8HM_VDC0#lF0qR5):tRRaAQ_Be a;m)R:YRRaAQ2CRs0MksRaQh )t ;R
R-)-RCD#k0kR#Lb0$CQ:Rhta  R)
RR--)kC#DR0:w8HM#ER0CCRDVF0l#F0ROsOksOCMCVRFRC0ERDPNkFCRVRRYHqMR)
t3R-R-RRRRRRRRR0)Ck#sMRC0ER8HMCFGRVER0CORFOsksCCMORRHVHC0RG0H##F,Rs4R-REF0CHsI#
C3
-RR-8RQ:3RqcR4
RMVkOF0HMHRVMs8_H0oEl0F#R)5qtRR:A_Qaea BmR);YRR:A2QaR0sCkRsMQ hat; )
-RR-CR)#0kDRL#k0C$b:hRQa  t)R
R-)-RCD#k0w:RH#M8RC0ERVDC0#lF0ORFOsksCCMORRFV0RECPkNDCVRFRHYRM)RqtR3
RR--RRRRRRRR)kC0sRM#0RECHCM8GVRFRC0EROFOkCssMROCHHVR0GRCH##0,sRFRR-4FC0Es#IHC
3
R-R-============================================================================
-RR-FRBlsbNHM#FRCmbsFN0sR#
R=--=========================================================================
==R-R-R:Q8R4B3
VRRk0MOHRFM"R>"5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B
3dRkRVMHO0F"MR>5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB6R
RVOkM0MHFR"">RR5p:QRAa _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNM-FMMNCo0CHPRaQh )t 3R

R=--=========================================================================
==R-R-R:Q8R(B3
VRRk0MOHRFM"R<"5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B
3gRkRVMHO0F"MR<5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB4R4
RMVkOF0HM<R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMF-oMCNP0HChRQa  t)
3
R-R-============================================================================
-RR-8RQ:3RB4Rd
RMVkOF0HM<R"=5"Rp),RRA:RQea_ mBa)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B634
VRRk0MOHRFM""<=RR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRHpR#RRNM-FMMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8R4B3(R
RVOkM0MHFR="<"pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMC-MoHN0PQCRhta  
)3
-RR-============================================================================R
R-Q-R8B:R3
4gRkRVMHO0F"MR>R="5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R.B34R
RVOkM0MHFR=">"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB.Rd
RMVkOF0HM>R"=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-=-==========================================================================R=
RR--QR8:B63.
VRRk0MOHRFM"R="5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B(3.
VRRk0MOHRFM"R="5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NFRMMC-MoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
.gRkRVMHO0F"MR=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"=pRRR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMC-MoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:B43d
VRRk0MOHRFM""/=R,5pR:)RRaAQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBdRd
RMVkOF0HM/R"=5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRRRH#NFRMMC-MoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
d6RkRVMHO0F"MR/R="5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNM-FMMNCo0CHPRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RBdR(
RMVkOF0HMQRvhzQvvpR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:QRAa _eB)am
-RR-CR)#0kD:CR)0Mks#ER0CCRD#s#CRRFV0RIFzQh1t7h ROPC0#FsRN0E0NRl$CRL
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBdRg
RMVkOF0HMQRvhzQvvpR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:A_Qaea BmR)
RR--)kC#DR0:)kC0sRM#0RECD#C#CFsRVRRNMMFMC0oNHRPCQ hat, )RRp,N
M8R-R-RRRRRRRRRRNMzQh1t7h ROPC0,FsR
)3
-RR-8RQ:3RBcR4
RMVkOF0HMQRvhzQvvpR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:A_Qaea BmR)
RR--)kC#DR0:)kC0sRM#0RECD#C#CFsRVMRNR1zhQ th7CRPOs0F,,RpR8NM
-RR-RRRRRRRRRRNMMFMC0oNHRPCQ hat, )R
)3
-RR-============================================================================R

RR--QR8:Bd3c
VRRk0MOHRFMvQqXvRzv5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:A_Qaea BmR)
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsF0VRIzFRht1QhR 7P0COFRs#00ENR$lNR
LCR-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RcB36R
RVOkM0MHFRXvqQvvzRR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CA:RQea_ mBa)R
R-)-RCD#k0):RCs0kM0#REoCRs0CNCFsRVRRNMMFMC0oNHRPCQ hat, )RRp,N
M8R-R-RRRRRRRRRRNMzQh1t7h ROPC0,FsR
)3
-RR-8RQ:3RBcR(
RMVkOF0HMqRvXzQvvpR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:A_Qaea BmR)
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsFNVRMhRz1hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRRMMFMNCo0CHPRaQh )t ,3R)
R
R-=-==========================================================================R=
RR--QR8:Bg3c
VRRk0MOHRFM""?>R,5pR:)RRaAQ_Be a2m)R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R6B34R
RVOkM0MHFR>"?"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:Bd36
VRRk0MOHRFM""?>RR5p:QRAa _eB)am;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R6B36R
RVOkM0MHFR<"?"pR5,RR):QRAa _eB)am2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB6R(
RMVkOF0HM?R"<5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RRMMFMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8R6B3gR
RVOkM0MHFR<"?"pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RBnR4
RMVkOF0HM?R"<R="5Rp,)RR:A_Qaea BmR)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RnB3dR
RVOkM0MHFR<"?=5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBnR6
RMVkOF0HM?R"<R="5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8RnB3(R
RVOkM0MHFR>"?=5"Rp),RRA:RQea_ mBa)s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bg3n
VRRk0MOHRFM"=?>"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRMMFMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8R(B34R
RVOkM0MHFR>"?=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:Bd3(
VRRk0MOHRFM""?=R,5pR:)RRaAQ_Be a2m)R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"=pRRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R(B36R
RVOkM0MHFR="?"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:B(3(
VRRk0MOHRFM""?=RR5p:QRAa _eB)am;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R(B3gR
RVOkM0MHFR/"?=5"Rp),RRA:RQea_ mBa)s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B43U
VRRk0MOHRFM"=?/"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RRMMFMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8RUB3dR
RVOkM0MHFR/"?=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R
R-1-RE0HVR8NMR0)FNR0CwOkM0MHF#R
R-=-==========================================================================
=
R-R-R:Q8R413
VRRk0MOHRFM1w]Qa _pw5aRqR)t:QRAa _eB)am;mRBzRha:qRhaqz)ps2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRussVFlN#RRH#EVD0-CRV0FNMRMhRz1hQt P7RCFO0smRBzRha0CHl#R3
RR--RRRRRRRRaRECPNNO0RC8bHF#0MHF#sRNCHRVD8DCR0IHEjR''R3
RR--RRRRRRRRaRECBhmzaCRDVF0l#C0RDCClMR0#NRsCD0F#3R

RR--QR8:1
3.RkRVMHO0F1MR]aQw_t)Q]5aRqR)t:QRAa _eB)am;mRBzRha:qRhaqz)ps2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slR#NRE0HV-osHEF0RMMRNR1zhQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0R''j3R
R-R-RRRRRRaRREBCRmazhRosHEF0l#C0RDCClMR0#NRsCD0F#3R
R-=-==========================================================================
=
R-R-R:Q8R613
VRRk0MOHRFM)qmaap _ Rwa5tq)RA:RQea_ mBa)B;RmazhRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFqs5)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NFRs0CN0-VDC0VRFRRNMzQh1t7h ROPC0RFsBhmzaHR0l3C#
R
R-Q-R81:R3Rn
RMVkOF0HMmR)a qa_t)Q]5aRqR)t:QRAa _eB)am;mRBzRha:qRhaqz)ps2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CL:RHP0_CFO0s)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRussVFlN#RR0sFN-0CsEHo0VRFRRNMzQh1t7h ROPC0RFsBhmzaHR0l3C#
R

R=--=========================================================================
==
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R1g#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R1gR
RVOkM0MHFRD"#D5"RqR)t:QRAa _eB)am;mRBzRha:hRQa  t)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CA:RQea_ mBa))5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:]R1Q_wapa w5tq),mRBz2ha
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0F1MR3R44HM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1434
VRRk0MOHRFM"D#s"qR5):tRRaAQ_Be a;m)RzBmh:aRRaQh )t 2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:QRAa _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]w)a_Qat]5tq),mRBz2ha
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0F1MR3R4dHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1d34
VRRk0MOHRFM"DsF"qR5):tRRaAQ_Be a;m)RzBmh:aRRaQh )t 2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:QRAa _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a pa w5tq),mRBz2ha
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0F1MR3R46HM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1634
VRRk0MOHRFM"ssF"qR5):tRRaAQ_Be a;m)RzBmh:aRRaQh )t 2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:QRAa _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a )]Qta)5qtB,Rmazh2R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1(34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413(R
RVOkM0MHFRD"#N5"RqR)t:QRAa _eB)am;mRBzRha:hRQa  t)s2RCs0kMQRAa _eB)am;R
R-)-RCD#k0kR#Lb0$CA:RQea_ mBa))5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:]R1Q_wapa w5tq),mRBz2ha
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0F1MR3R4gHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1g34
VRRk0MOHRFM"N#s"qR5):tRRaAQ_Be a;m)RzBmh:aRRaQh )t 2CRs0MksRaAQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:QRAa _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]w)a_Qat]5tq),mRBz2ha
R

R=--=========================================================================
==R-R-R)RR Z1Q kRwMHO0F
M#R-R-============================================================================
R
R-Q-R8):R3R.
RMVkOF0HM R)1 QZR)5qtRR:A_Qaea BmR);h_ W1 QZRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COFhs5 1W_Q-Z 4FR8IFM0R
j2R-R-R#)Ck:D0R#)CH#xCRC0ER1zhQ th7CRPOs0FRtq)RR0F0REC#ObCHCVH8HR#x
C3R-R-RRRRRRRRRRaFONsC0NCRRsDNoRCsP0COFRs,0RECMRCIrVDC0#lF0L9RHb0RF0#HH#FM
-RR-RRRRRRRRsRNCHRVD8DCR0IHEjR''W3RERCM0MskOHN0MRo,0RECD0CVl0F#R0LH#R
R-R-RRRRRRNRRs8CRsbFbC
83
VRRk0MOHRFM)Q 1Z5 Rq,)tRZ1Q  _)1RR:A_Qaea BmR)2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:A_Qaea Bm5)R1 QZ_1) 'MDCo-0E4FR8IFM0R
j2
-RR-============================================================================R
R-B-RFCMPsF#HMkRwMHO0F
M#R-R-============================================================================
R
R-Q-R87:R3R4
RMVkOF0HMmRa_aQh )t R)5qtRR:A_Qaea BmR)2skC0shMRq)azq
p;R-R-R#)CkRD0#0kL$:bCRahqzp)q3NReDRkCOMNMFL0RCCRMoHN0P#CRHCMORsbNN0lCCHsR#MRN
-RR-RRRRRRRRRRRRhRz1hQt P7RCFO0sR3
RR--)kC#DR0:BPFMC#s0RC0ER1zhQ th7CRPOs0FRR0FNQMRhta  
)3
-RR-8RQ:3R7dR
RVOkM0MHFR_aFAeH0CFO0sqR5)Rt,1 QZRh:Rq)azqRp2skC0sAMRQea_ mBa)R;
RR--)kC#D#0Rk$L0bRC:L_H0P0COF1s5Q-Z 4FR8IFM0R
j2R-R-R#)Ck:D0RMBFP0Cs#RRNM-FMMNCo0CHPRaQh )t RR0FNzMRht1QhR 7P0COFIsRH
0ER-R-RRRRRRRRRC0ERC#bOHHVC#8RH3xC
R
RVOkM0MHFR_aFAeH0CFO0sqR5):tRRahqzp)q;QR1Z) _ :1RRaAQ_Be a2m)
RRRR0sCkRsMA_Qaea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_tpmQeB_ mBa)Q51Z) _ D1'C0MoER-48MFI0jFR2-

-CRLoRHMp-B1.njj-j4d
NRRD#HNR_aFA_H0e0COFHsR#R
RRFRa_0AHe0COFhsrq)azqRp,hzqa)RqpskC0sAMRQea_ mBa)
9;RDRNHRN#aAF_e#RH
RRRR_aFAeH0CFO0sqrhaqz)ph,Rq)azqspRCs0kMQRAa _eB)am9
;
RDRNHRN#aAF_He0_CFO0s#RH
RRRR_aFAeH0CFO0sqrhaqz)pA,RQea_ mBa)CRs0MksRaAQ_Be a9m);R
RNNDH#FRa_RAeHR#
RaRRFH_A0OeC0rFshzqa),qpRaAQ_Be aRm)skC0sAMRQea_ mBa)
9;
8CMRObN	CNoRvhz B)Q_aAQ_1zhQ th7
;
DsHLNRs$HCCC;#
kCCRHCMC3kslCHLO_HN03D
D;
ObN	CNoR8LF$zRhvQ )BQ_Aah_z1hQt H7R#R

RR--QR8:q
3dRkRVMHO0F"MR+5"Rp),RRA:RQea_ mBa)s2RCs0kMQRAa _eB)amR
H#RCRLo
HMRRRRskC0sAMRQea_ mBa)zR5ht1Qh5 7p+2RR1zhQ th725)2R;
R8CMRMVkOF0HM+R""
;
R-R-R:Q8Rdq3)R
RVOkM0MHFR""+5:pRRaAQ_Be a;m)R:)RRaAQ2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt p752RR+)
2;RMRC8kRVMHO0F"MR+
";
-RR-8RQ:3RqdRp
RMVkOF0HM+R""R5p:QRAa);RRA:RQea_ mBa)s2RCs0kMQRAa _eB)amR
H#RCRLo
HMRRRRskC0sAMRQea_ mBa)pR5Rz+Rht1Qh5 7);22
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3R6
RMVkOF0HM+R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2+2R);R
RCRM8VOkM0MHFR""+;R

RR--QR8:q
3nRkRVMHO0F"MR+5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)5+pRR1zhQ th725)2R;
R8CMRMVkOF0HM+R""
;
R-R-============================================================================
R
R-Q-R8q:R3Rg
RMVkOF0HM-R""pR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt p752RR-zQh1t7h 52)2;R
RCRM8VOkM0MHFR""-;R

RR--QR8:q)3g
VRRk0MOHRFM"5-"pRR:A_Qaea BmR);)RR:A2QaR0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)51zhQ th725pR)-R2R;
R8CMRMVkOF0HM-R""
;
R-R-R:Q8Rgq3pR
RVOkM0MHFR""-5:pRRaAQ;RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRR5p-hRz1hQt )752
2;RMRC8kRVMHO0F"MR-
";
-RR-8RQ:3Rq4R4
RMVkOF0HM-R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2-2R);R
RCRM8VOkM0MHFR""-;R

RR--QR8:q.34
VRRk0MOHRFM"R-"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRR5p-hRz1hQt )752
2;RMRC8kRVMHO0F"MR-
";
-RR-============================================================================R

RR--QR8:q634
VRRk0MOHRFM"R*"5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2*hRz1hQt )752
2;RMRC8kRVMHO0F"MR*
";
-RR-8RQ:3Rq4R(
RMVkOF0HM*R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2*2R);R
RCRM8VOkM0MHFR""*;R

RR--QR8:qU34
VRRk0MOHRFM"R*"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRR5p*hRz1hQt )752
2;RMRC8kRVMHO0F"MR*
";
-RR-============================================================================R

RR--QR8:q43.
VRRk0MOHRFM"R/"5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2/hRz1hQt )752
2;RMRC8kRVMHO0F"MR/
";
-RR-8RQ:3Rq.Rd
RMVkOF0HM/R""pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2/2R);R
RCRM8VOkM0MHFR""/;R

RR--QR8:qc3.
VRRk0MOHRFM"R/"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRR5p/hRz1hQt )752
2;RMRC8kRVMHO0F"MR/
";
-RR-============================================================================R

RR--QR8:q(3.
VRRk0MOHRFM"lsC"pR5,RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt p752CRslhRz1hQt )752
2;RMRC8kRVMHO0F"MRs"Cl;R

RR--QR8:qg3.
VRRk0MOHRFM"lsC"pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2sRCl)
2;RMRC8kRVMHO0F"MRs"Cl;R

RR--QR8:qj3d
VRRk0MOHRFM"lsC"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RpCRslhRz1hQt )752
2;RMRC8kRVMHO0F"MRs"Cl;R

R=--=========================================================================
==
-RR-8RQ:3RqdRd
RMVkOF0HMlR"FR8"5Rp,)RR:A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5Rp2lRF8zQh1t7h 52)2;R
RCRM8VOkM0MHFRF"l8
";
-RR-8RQ:3RqdR6
RMVkOF0HMlR"FR8"5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt p752FRl82R);R
RCRM8VOkM0MHFRF"l8
";
-RR-8RQ:3RqdRn
RMVkOF0HMlR"FR8"5:pRRahqzp)q;RR):QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRR5plRF8zQh1t7h 52)2;R
RCRM8VOkM0MHFRF"l8
";
-RR-============================================================================R
R-Q-R8q:R3
dgRkRVMHO0FVMRH_M8D0CVl0F#R)5qtA:RQea_ mBa)Y;R:QRAas2RCs0kMhRQa  t)#RH
LRRCMoH
RRRR0sCkRsMV8HM_VDC0#lF0h5z1hQt q75),t2R;Y2
CRRMV8Rk0MOHRFMV8HM_VDC0#lF0
;
R-R-R:Q8Rcq34R
RVOkM0MHFRMVH8H_solE0FR#05tq):QRAa _eB)am;:RYRaAQ2CRs0MksRaQh )t R
H#RCRLo
HMRRRRskC0sVMRH_M8sEHo0#lF0h5z1hQt q75),t2R;Y2
CRRMV8Rk0MOHRFMV8HM_osHEF0l#
0;
-RR-============================================================================R
R-Q-R8B:R3R4
RMVkOF0HM>R""pR5,RR):QRAa _eB)am2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p>2RR1zhQ th725);R
RCRM8VOkM0MHFR"">;R

RR--QR8:B
3dRkRVMHO0F"MR>5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMRRp>hRz1hQt )752R;
R8CMRMVkOF0HM>R""
;
R-R-R:Q8R6B3
VRRk0MOHRFM"R>"5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p>2RR
);RMRC8kRVMHO0F"MR>
";
-RR-============================================================================R
R-Q-R8B:R3R(
RMVkOF0HM<R""pR5,RR):QRAa _eB)am2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p<2RR1zhQ th725);R
RCRM8VOkM0MHFR""<;R

RR--QR8:B
3gRkRVMHO0F"MR<5"RpRR:hzqa);qpR:)RRaAQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMRRp<hRz1hQt )752R;
R8CMRMVkOF0HM<R""
;
R-R-R:Q8R4B34R
RVOkM0MHFR""<RR5p:QRAa _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2<;R)
CRRMV8Rk0MOHRFM";<"
R
R-=-==========================================================================R=
RR--QR8:Bd34
VRRk0MOHRFM""<=R,5pR:)RRaAQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752=R<R1zhQ th725);R
RCRM8VOkM0MHFR="<"
;
R-R-R:Q8R4B36R
RVOkM0MHFR="<"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR<pR=hRz1hQt )752R;
R8CMRMVkOF0HM<R"=
";
-RR-8RQ:3RB4R(
RMVkOF0HM<R"=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752=R<R
);RMRC8kRVMHO0F"MR<;="
R
R-=-==========================================================================R=
RR--QR8:Bg34
VRRk0MOHRFM"">=R,5pR:)RRaAQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752=R>R1zhQ th725);R
RCRM8VOkM0MHFR=">"
;
R-R-R:Q8R.B34R
RVOkM0MHFR=">"pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR>pR=hRz1hQt )752R;
R8CMRMVkOF0HM>R"=
";
-RR-8RQ:3RB.Rd
RMVkOF0HM>R"=5"RpRR:A_Qaea BmR);)RR:hzqa)2qpR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752=R>R
);RMRC8kRVMHO0F"MR>;="
R
R-=-==========================================================================R=
RR--QR8:B63.
VRRk0MOHRFM"R="5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRz=Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR=
";
-RR-8RQ:3RB.R(
RMVkOF0HM=R""pR5Rh:Rq)azqRp;)RR:A_Qaea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR=pRR1zhQ th725);R
RCRM8VOkM0MHFR""=;R

RR--QR8:Bg3.
VRRk0MOHRFM"R="5:pRRaAQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p=2RR
);RMRC8kRVMHO0F"MR=
";
-RR-============================================================================R
R-Q-R8B:R3
d4RkRVMHO0F"MR/R="5Rp,)RR:A_Qaea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR/=zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""/=;R

RR--QR8:Bd3d
VRRk0MOHRFM""/=RR5p:qRhaqz)p);RRA:RQea_ mBa)s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMp=R/R1zhQ th725);R
RCRM8VOkM0MHFR="/"
;
R-R-R:Q8RdB36R
RVOkM0MHFR="/"pR5RA:RQea_ mBa));RRh:Rq)azqRp2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR/=)R;
R8CMRMVkOF0HM/R"=
";
-RR-============================================================================R
R-Q-R8B:R3
d(RkRVMHO0FvMRQvhQz5vRp),R:QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRQ5vhzQvvh5z1hQt p752z,Rht1Qh5 7)222;R
RCRM8VOkM0MHFRhvQQvvz;R

RR--QR8:Bg3d
VRRk0MOHRFMvQQhvRzv5Rp:hzqa);qpRR):A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RvQQhv5zvpz,Rht1Qh5 7)222;R
RCRM8VOkM0MHFRhvQQvvz;R

RR--QR8:B43c
VRRk0MOHRFMvQQhvRzv5Rp:A_Qaea BmR);)h:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RvQQhv5zvzQh1t7h 5,p2R2)2;R
RCRM8VOkM0MHFRhvQQvvz;R

R=--=========================================================================
==R-R-R:Q8RcB3dR
RVOkM0MHFRXvqQvvzR,5pRR):A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RvQqXv5zvzQh1t7h 5,p2R1zhQ th725)2
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcR6
RMVkOF0HMqRvXzQvvpR5:qRhaqz)p);R:QRAa _eB)am2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRq5vXzQvv,5pR1zhQ th725)2
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcR(
RMVkOF0HMqRvXzQvvpR5:QRAa _eB)am;:R)Rahqzp)q2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRq5vXzQvvh5z1hQt p752),R2
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-============================================================================R

RR--QR8:Bg3c
VRRk0MOHRFM""?>R,5pRR):A_Qaea BmR)2skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?>zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:B436
VRRk0MOHRFM""?>R:5pRahqzp)q;:R)RaAQ_Be a2m)R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMRRp?z>Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR?;>"
R
R-Q-R8B:R3
6dRkRVMHO0F"MR?R>"5Rp:A_Qaea BmR);)h:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?>)R;
R8CMRMVkOF0HM?R">
";
-RR-============================================================================R

RR--QR8:B636
VRRk0MOHRFM""?<R,5pRR):A_Qaea BmR)2skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?<zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""?<;R

RR--QR8:B(36
VRRk0MOHRFM""?<R:5pRahqzp)q;:R)RaAQ_Be a2m)R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMRRp?z<Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
6gRkRVMHO0F"MR?R<"5Rp:A_Qaea BmR);)h:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?<)R;
R8CMRMVkOF0HM?R"<
";
-RR-============================================================================R

RR--QR8:B43n
VRRk0MOHRFM"=?<"pR5,:R)RaAQ_Be a2m)R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752<R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
ndRkRVMHO0F"MR?"<=R:5pRahqzp)q;:R)RaAQ_Be a2m)R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMRRp?R<=zQh1t7h 5;)2
CRRMV8Rk0MOHRFM"=?<"
;
R-R-R:Q8RnB36R
RVOkM0MHFR<"?=5"RpA:RQea_ mBa));R:qRhaqz)ps2RCs0kMQRAa#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2?R<=)R;
R8CMRMVkOF0HM?R"<;="
R
R-=-==========================================================================
=
R-R-R:Q8RnB3(R
RVOkM0MHFR>"?=5"Rp),R:QRAa _eB)am2CRs0MksRaAQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R>z=Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR?">=;R

RR--QR8:Bg3n
VRRk0MOHRFM"=?>"pR5:qRhaqz)p);R:QRAa _eB)am2CRs0MksRaAQR
H#RCRLo
HMRRRRskC0spMRR=?>R1zhQ th725);R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RB(R4
RMVkOF0HM?R">R="5Rp:A_Qaea BmR);)h:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR1zhQ th725pR=?>R
);RMRC8kRVMHO0F"MR?">=;R

R=--=========================================================================
==
-RR-8RQ:3RB(Rd
RMVkOF0HM?R"=5"Rp),R:QRAa _eB)am2CRs0MksRaAQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R=hRz1hQt )752R;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(R6
RMVkOF0HM?R"=5"Rph:Rq)azqRp;)A:RQea_ mBa)s2RCs0kMQRAa#RH
LRRCMoH
RRRR0sCkRsMp=R?R1zhQ th725);R
RCRM8VOkM0MHFR="?"
;
R-R-R:Q8R(B3(R
RVOkM0MHFR="?"pR5:QRAa _eB)am;:R)Rahqzp)q2CRs0MksRaAQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R=;R)
CRRMV8Rk0MOHRFM""?=;R

R=--=========================================================================
==
-RR-8RQ:3RB(Rg
RMVkOF0HM?R"/R="5Rp,)A:RQea_ mBa)s2RCs0kMQRAa#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2?R/=zQh1t7h 5;)2
CRRMV8Rk0MOHRFM"=?/"
;
R-R-R:Q8RUB34R
RVOkM0MHFR/"?=5"Rph:Rq)azqRp;)A:RQea_ mBa)s2RCs0kMQRAa#RH
LRRCMoH
RRRR0sCkRsMp/R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"/;="
R
R-Q-R8B:R3
UdRkRVMHO0F"MR?"/=R:5pRaAQ_Be a;m)RR):hzqa)2qpR0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752/R?=;R)
CRRMV8Rk0MOHRFM"=?/"
;
R-R-============================================================================
R
R-Q-R81:R3R4
RMVkOF0HM]R1Q_wapa wR)5qtRR:A_Qaea BmR);BhmzaRR:hzqa)2qpR0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)5H#EVD0_CRV05tq)R=RR>hRz1hQt q75),t2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBhmza>R=RzBmh2a2;R
RCRM8VOkM0MHFRQ1]wpa_ ;wa
R
R-Q-R81:R3R.
RMVkOF0HM]R1Q_wa)]QtaqR5):tRRaAQ_Be a;m)RzBmh:aRRahqzp)q2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRE5#H_V0sEHo0qR5)RtRRR=>zQh1t7h 5tq)2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBRRmazhRR=>Bhmza;22
CRRMV8Rk0MOHRFM1w]QaQ_)t;]a
R
R-=-==========================================================================
=
R-R-R:Q8R613
VRRk0MOHRFM)qmaap _ Rwa5tq)RA:RQea_ mBa)B;RmazhRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RsNF00DC_CRV05tq)R=RR>hRz1hQt q75),t2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRzBmh=aR>mRBz2ha2R;
R8CMRMVkOF0HMmR)a qa_wp a
;
R-R-R:Q8Rn13
VRRk0MOHRFM)qmaa) _Qat]R)5qtRR:A_Qaea BmR);BhmzaRR:hzqa)2qpR0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)50sFN_0CsEHo0qR5)RtRRR=>zQh1t7h 5tq)2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRBhmza>R=RzBmh2a2;R
RCRM8VOkM0MHFRa)mq_a )]Qta
;
R-R-============================================================================
R
R-Q-R81:R3Rg
RMVkOF0HM#R"DRD"5tq):QRAa _eB)am;mRBz:haRaQh )t 2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt q75)Rt2#RDDBhmza
2;RMRC8kRVMHO0F"MR#"DD;R

RR--QR8:1434
VRRk0MOHRFM"D#s"qR5)Rt:A_Qaea BmR);BhmzaQ:Rhta  R)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5tq)2sR#DmRBz2ha;R
RCRM8VOkM0MHFRs"#D
";
-RR-8RQ:3R14Rd
RMVkOF0HMsR"FRD"5tq):QRAa _eB)am;mRBz:haRaQh )t 2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt q75)Rt2sRFDBhmza
2;RMRC8kRVMHO0F"MRs"FD;R

RR--QR8:1634
VRRk0MOHRFM"ssF"qR5)Rt:A_Qaea BmR);BhmzaQ:Rhta  R)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5tq)2FRssmRBz2ha;R
RCRM8VOkM0MHFRF"ss
";
-RR-8RQ:3R14R(
RMVkOF0HM#R"DRN"5tq):QRAa _eB)am;mRBz:haRaQh )t 2CRs0MksRaAQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMQRAa _eB)amRh5z1hQt q75)Rt2#RDNBhmza
2;RMRC8kRVMHO0F"MR#"DN;R

RR--QR8:1g34
VRRk0MOHRFM"N#s"qR5)Rt:A_Qaea BmR);BhmzaQ:Rhta  R)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)RzQh1t7h 5tq)2sR#NmRBz2ha;R
RCRM8VOkM0MHFRs"#N
";
-RR-============================================================================R

RR--QR8:)
3.RkRVMHO0F)MR Z1Q qR5):tRRaAQ_Be a;m)RWh _Z1Q RR:hzqa)2qpR0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)5R
RRRRRsHC#x5CRNRsoRRRRRR=>zQh1t7h 5tq)2R,
RRRRRRRRRRRRRWh _Z1Q >R=RWh _Z1Q ;22
CRRMV8Rk0MOHRFM)Q 1Z
 ;
VRRk0MOHRFM)Q 1Z5 Rq,)tRZ1Q  _)1RR:A_Qaea BmR)2skC0sAMRQea_ mBa)#RH
LRRCMoH
RRRR0sCkRsMA_Qaea Bm5)R
RRRR)RR Z1Q qR5)RtRRRRR=z>Rht1Qh5 7q2)t,R
RRRRRRRRRRRRRh_ W1 QZRR=>1 QZ_1) 'MDCo20E2R;
R8CMRMVkOF0HM R)1 QZ;R

R=--=========================================================================
==
-RR-8RQ:3R74R
RVOkM0MHFR_amQ hatR )5tq)RA:RQea_ mBa)s2RCs0kMqRhaqz)p#RH
LRRCMoH
RRRR0sCkRsMaQm_hta  5)RzQh1t7h 5tq)2
2;RMRC8kRVMHO0FaMRmh_Qa  t)
;
R-R-R:Q8Rd73
VRRk0MOHRFMaAF_HC0eOs0FR)5qt1,RQRZ :qRhaqz)ps2RCs0kMQRAa _eB)amR
H#RCRLo
HMRRRRskC0sAMRQea_ mBa)aR5mh_z1hQt q75)Rt,1 QZ2
2;RMRC8kRVMHO0FaMRFH_A0OeC0;Fs
R
RVOkM0MHFR_aFAeH0CFO0sqR5):tRRahqzp)q;QR1Z) _ :1RRaAQ_Be a2m)
RRRR0sCkRsMA_Qaea BmH)R#R
RLHCoMR
RRCRs0MksRaAQ_Be aRm)5_amzQh1t7h 5tq),QR1Z) _ D1'C0MoE;22
CRRMV8Rk0MOHRFMaAF_HC0eOs0F;C

Mb8RNNO	oLCRFR8$h zv)_QBA_QazQh1t7h ;



