--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb/oIlbNbC/s#GHHDMDG/HoL/CsMCHoO/CoM_CsMCH/O.s_Nls3IbPyE84
Rf-
-
---
--
-Rl1HbRDC)RqvIEH0RM#HoRDCq)77 R11VRFsLEF0RNsC8MRN8sRIH
0C-a-RNCso0RR:XHHDM-G
-D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
0CMHR0$)_qv)RWuHS#
oCCMsRHO5S
SVHNlD:$RRs#0HRMo:"=RMCFM"S;
S8IH0:ERR0HMCsoCRR:=.
;RS8SN8HsI8R0E:MRH0CCos=R:RRU;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0SE
Sb8C0:ERR0HMCsoCRR:=.;6n
8SSF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoS
S8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCSo
S8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRR-R-R8ENR8N8s#C#RosC
2SS;b
SFRs05S
S7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
S7RQhRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
Sq)77RH:RM0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;S
SWR R:MRHR8#0_oDFHRO;RRRRR-R-RHIs0CCRMDNLCFRVsNRslS
SBRpi:MRHR8#0_oDFHRO;RRRRR-R-RFODOV	RFssRNRl,Ns88,HR8MS
SmiBpRH:RM0R#8F_DoRHORRRRR-R-R0FbRFODOV	RF8sRF
k0S;S2
8CMR0CMHR0$)_qv);Wu
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCDRLF_O	sRNlF)VRq)v_WHuR#$
0bHCRMN0_s$sNRRH#NNss$jR5RR0F6F2RVMRH0CCosO;
F0M#NRM0I0H8Es_NsRN$:MRH0s_NsRN$:5=R4.,R,,RcRRg,4RU,d;n2
MOF#M0N0CR8b_0ENNss$RR:H_M0NNss$=R:Rn54d,UcRgU4.c,Rj,gnRc.jU4,Rj,.cR.642O;
F0M#NRM08dHP.RR:HCM0oRCs:5=RI0H8E2-4/;dn
MOF#M0N0HR8PR4n:MRH0CCos=R:RH5I8-0E442/UO;
F0M#NRM08UHPRH:RMo0CC:sR=IR5HE80-/42gO;
F0M#NRM08cHPRH:RMo0CC:sR=IR5HE80-/42cO;
F0M#NRM08.HPRH:RMo0CC:sR=IR5HE80-/42.O;
F0M#NRM084HPRH:RMo0CC:sR=IR5HE80-/424
;
O#FM00NMRFLFD:4RRFLFDMCNRR:=5P8H4RR>j
2;O#FM00NMRFLFD:.RRFLFDMCNRR:=5P8H.RR>j
2;O#FM00NMRFLFD:cRRFLFDMCNRR:=5P8HcRR>j
2;O#FM00NMRFLFD:URRFLFDMCNRR:=5P8HURR>j
2;O#FM00NMRFLFDR4n:FRLFNDCM=R:RH58PR4n>2Rj;F
OMN#0ML0RFdFD.RR:LDFFCRNM:5=R8dHP.RR>j
2;
MOF#M0N0HR8Pd4nU:cRR0HMCsoCRR:=5b8C04E-2n/4d;Uc
MOF#M0N0HR8PgU4.RR:HCM0oRCs:5=R80CbE2-4/gU4.O;
F0M#NRM08cHPjRgn:MRH0CCos=R:RC58b-0E4c2/j;gn
MOF#M0N0HR8Pc.jURR:HCM0oRCs:5=R80CbE2-4/c.jUO;
F0M#NRM084HPjR.c:MRH0CCos=R:RC58b-0E442/j;.c
MOF#M0N0HR8P.64RH:RMo0CC:sR=8R5CEb0-/426;4.
F
OMN#0ML0RF6FD4:.RRFLFDMCNRR:=5P8H6R4.>2Rj;F
OMN#0ML0RF4FDjR.c:FRLFNDCM=R:RH58P.4jcRR>j
2;O#FM00NMRFLFDc.jURR:LDFFCRNM:5=R8.HPjRcU>2Rj;F
OMN#0ML0RFcFDjRgn:FRLFNDCM=R:RH58PgcjnRR>j
2;O#FM00NMRFLFDgU4.RR:LDFFCRNM:5=R8UHP4Rg.>2Rj;F
OMN#0ML0RF4FDncdURL:RFCFDN:MR=8R5HnP4dRUc>2Rj;O

F0M#NRM0#_klI0H8ERR:HCM0oRCs:A=Rm mpqbh'FL#5F4FD2RR+Apmm 'qhb5F#LDFF.+2RRmAmph q'#bF5FLFDRc2+mRAmqp hF'b#F5LF2DURA+Rm mpqbh'FL#5F4FDn
2;O#FM00NMRl#k_b8C0:ERR0HMCsoCRR:=6RR-5mAmph q'#bF5FLFD.642RR+Apmm 'qhb5F#LDFF4cj.2RR+Apmm 'qhb5F#LDFF.Ujc2RR+Apmm 'qhb5F#LDFFcnjg2RR+Apmm 'qhb5F#LDFFU.4g2
2;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lH_I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5kIl_HE802O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_kl80CbE
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_b8C0;E2
F
OMN#0MI0R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/42IE_OFCHO_8IH0+ERR
4;O#FM00NMR8I_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/IOHEFO8C_CEb0R4+R;O

F0M#NRM08H_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/O8_EOFHCH_I8R0E+;R4
MOF#M0N0_R880CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E482/_FOEH_OC80CbERR+4
;
O#FM00NMR#I_HRxC:MRH0CCos=R:RII_HE80_lMk_DOCD*#RR8I_CEb0_lMk_DOCD
#;O#FM00NMR#8_HRxC:MRH0CCos=R:RI8_HE80_lMk_DOCD*#RR88_CEb0_lMk_DOCD
#;
MOF#M0N0FRLF8D_RL:RFCFDN:MR=8R5_x#HCRR-IH_#x<CR=2Rj;F
OMN#0ML0RF_FDIRR:LDFFCRNM:M=RFL05F_FD8
2;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_8IH0;E2
MOF#M0N0EROFCHO_b8C0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_b8C0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*H5I8-0E482/_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*80CbE2-4/O8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4
O--F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8R-F-OMN#0MD0RC_V0FsPCRH:RMo0CC:sR=5R55b8C0+ERR246R8lFR2d.R4/RnR2;RRRRRRRRRRRRRRRRRRRRRRRR-y-RRRFV)4qvn1X4RCMC8RC8VRFsD0CVRCFPsFRIs
8#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD8RNsRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-R-RR0FsHCo#s0CRC0ERD#CCRO0#MHoNFDRVsR0HN#00NC
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjj"RR&Ns8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj&"RR_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjRj"&8RN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjj"jjRN&R8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FINs88RR<="jjjj&"RR_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FINs88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R''jRN&R8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FINs88RR<=Ns8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR4RnR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRR(z4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4(
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRp-i
-RRRRnz4RRR:H5VRNs88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCH-M
-RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Cz;4n
R--RzRR4:(RRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);-C-SMo8RCsMCNR0Cz;4(
RSRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>cR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRc<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;c2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.j:VRHR85N8HsI8R0E>cR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4RR:)Aqv41n_4R
SRRRRRRRRRbRRFRs0lRNb557Qj=2R>MRH_osC5,[2R7q7)>R=RIDF_8N8sd54RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57mj=2R>kRF0k_L#H45,2[2;R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRSRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>dR42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFdR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRd
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.RX.:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvU.4gX:.RRv)qA_4n1S.
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7=)R>FRDI8_N84s5.FR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R42=F>RkL0_k5#.H*,.[2+4,mR75Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR.<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;.2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnXRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gcjnRXc:qR)vnA4_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7R7)=D>RFNI_858s484RF0IMF2Rj,hR RR=>',4'R)11RR=>',j'RS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25dRR=>F_k0Lck#5RH,c+*[dR2,7.m52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSS57m4=2R>kRF0k_L#Hc5,[c*+,42R57mj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1
dSzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>R4o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR4<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;42
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUXRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_c.jURXU:qR)vnA4_
1gSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7R7)=D>RFNI_858s48jRF0IMF2Rj,hR RR=>',4'R)11RR=>',j'RS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25(RR=>F_k0LUk#5UH,*([+27,Rm25nRR=>F_k0LUk#5UH,*n[+2
,RSSSS76m52>R=R0Fk_#LkU,5HU+*[6R2,7cm52>R=R0Fk_#LkU,5HU+*[cR2,7dm52>R=R0Fk_#LkU,5HU+*[dR2,
SSSS57m.=2R>kRF0k_L#HU5,[U*+,.2R57m4=2R>kRF0k_L#HU5,[U*+,42R57mj=2R>kRF0k_L#HU5,[U*2
,RSSSS75Quj=2R>MRH_osC5[g*+,U2Ru7m5Rj2=b>RN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH[,R2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>RjRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rj2<N=R8C_so85N8HsI8-0E4FR8IFM0R24j;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;cj
-S-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRcSz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;c4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4:nRRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_jX.c4:nRRv)qA_4n1
4USRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7=)R>FRDI8_N8gs5RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4R62=F>RkL0_kn#454H,n+*[4,62R57m4Rc2=F>RkL0_kn#454H,n+*[4,c2RS
SSmS7524dRR=>F_k0L4k#n,5H4[n*+24d,mR7524.RR=>F_k0L4k#n,5H4[n*+24.,mR75244RR=>F_k0L4k#n,5H4[n*+244,SR
S7SSmj542>R=R0Fk_#Lk4Hn5,*4n[j+427,Rm25gRR=>F_k0L4k#n,5H4[n*+,g2R57mU=2R>kRF0k_L#54nHn,4*U[+2S,
S7SSm25(RR=>F_k0L4k#n,5H4[n*+,(2R57mn=2R>kRF0k_L#54nHn,4*n[+27,Rm256RR=>F_k0L4k#n,5H4[n*+,62
SSSRRRR7cm52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR75Rd2=F>RkL0_kn#454H,n+*[dR2,7.m52>R=R0Fk_#Lk4Hn5,*4n[2+.,S
SRRRRRRRR74m52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR75Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+n
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_kn#45RH,.+*[4R2,75muj=2R>NRbs$H0_#Lk4Hn5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRc
.;RRRRRMSC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nz
Sc:dRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR2gRRMoCC0sNCR
SRzRRO:D	RFbsO#C#Rp5BiS2
SLRRCMoH
RSSRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRSRRRRRNC8so85N8HsI8-0E4FR8IFM0RRg2<N=R8C_so85N8HsI8-0E4FR8IFM0R;g2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;SRRRRczcRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SS6zcRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SFSSkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc
6;SR--Q5VRNs88I0H8E=R<RRg2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
SSSzRcn:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzRc(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRR)RAq6v_4d.X.RR:)Aqv41n_dRn
RRRRRRRRRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77RD=>FNI_858sUFR8IFM0R,j2RR h='>R4R',1R1)='>Rj
',RRRRRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm45d2>R=R0Fk_#LkdH.5,*d.[4+d27,Rmj5d2>R=R0Fk_#LkdH.5,*d.[j+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rg2=F>RkL0_k.#d5dH,.+*[.,g2R57m.RU2=F>RkL0_k.#d5dH,.+*[.,U2R57m.R(2=F>RkL0_k.#d5dH,.+*[.,(2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmn5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rmc5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rd2=F>RkL0_k.#d5dH,.+*[.,d2R57m.R.2=F>RkL0_k.#d5dH,.+*[.,.2R57m.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rmg542>R=R0Fk_#LkdH.5,*d.[g+427,RmU542>R=R0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4R(2=F>RkL0_k.#d5dH,.+*[4,(2R57m4Rn2=F>RkL0_k.#d5dH,.+*[4,n2R57m4R62=F>RkL0_k.#d5dH,.+*[4,62
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmc542>R=R0Fk_#LkdH.5,*d.[c+427,Rmd542>R=R0Fk_#LkdH.5,*d.[d+427,Rm.542>R=R0Fk_#LkdH.5,*d.[.+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75244RR=>F_k0Ldk#.,5Hd[.*+244,mR7524jRR=>F_k0Ldk#.,5Hd[.*+24j,mR75Rg2=F>RkL0_k.#d5dH,.+*[gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm25URR=>F_k0Ldk#.,5Hd[.*+,U2R57m(=2R>kRF0k_L#5d.H.,d*([+27,Rm25nRR=>F_k0Ldk#.,5Hd[.*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR76m52>R=R0Fk_#LkdH.5,*d.[2+6,mR75Rc2=F>RkL0_k.#d5dH,.+*[cR2,7dm52>R=R0Fk_#LkdH.5,*d.[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.=2R>kRF0k_L#5d.H.,d*.[+27,Rm254RR=>F_k0Ldk#.,5Hd[.*+,42R57mj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,Rmdu52>R=RsbNH_0$Ldk#.,5HR[c*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.u52>R=RsbNH_0$Ldk#.,5HR[c*+,.2Ru7m5R42=b>RN0sH$k_L#5d.Hc,R*4[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5Rj2=b>RN0sH$k_L#5d.Hc,R*2[2;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SCSSMo8RCsMCNR0Cz;c(
CSSMo8RCsMCNR0Cz;cc
MSC8CRoMNCs0zCRc
d;CRM8NEsOHO0C0CksRFLDOs	_N
l;
R--MsF_IE_OCRO	VRFs#oHMDbCRFRs0)RqvHH#R80CMHDONRR0FLODF	NRsls
NO0EHCkO0sMCRFI_s_COEOF	RVqR)vW_)u#RH
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVMsF_IE_OCRO	:sRNO0EHCkO0sHCR#zR"#oHMRFLDOs	_NVlRF#sRHDMoCFRbss0RNIlRHR0E#_$Ms#Nl0C$DR_MFsOI_E	CO"0;
$RbCH_M0NNss$#RHRsNsN5$RjFR0RR62FHVRMo0CC
s;O#FM00NMR8IH0NE_s$sNRH:RMN0_s$sNRR:=5R4,.c,R,,RgR,4UR2dn;F
OMN#0M80RCEb0_sNsN:$RR0HM_sNsN:$R=4R5ncdU,4RUgR.,cnjg,jR.cRU,4cj.,4R6.
2;O#FM00NMRP8Hd:.RR0HMCsoCRR:=58IH04E-2n/d;F
OMN#0M80RHnP4RH:RMo0CC:sR=IR5HE80-/424
U;O#FM00NMRP8HURR:HCM0oRCs:5=RI0H8E2-4/
g;O#FM00NMRP8HcRR:HCM0oRCs:5=RI0H8E2-4/
c;O#FM00NMRP8H.RR:HCM0oRCs:5=RI0H8E2-4/
.;O#FM00NMRP8H4RR:HCM0oRCs:5=RI0H8E2-4/
4;
MOF#M0N0FRLFRD4:FRLFNDCM=R:RH58P>4RR;j2
MOF#M0N0FRLFRD.:FRLFNDCM=R:RH58P>.RR;j2
MOF#M0N0FRLFRDc:FRLFNDCM=R:RH58P>cRR;j2
MOF#M0N0FRLFRDU:FRLFNDCM=R:RH58P>URR;j2
MOF#M0N0FRLFnD4RL:RFCFDN:MR=8R5HnP4Rj>R2O;
F0M#NRM0LDFFd:.RRFLFDMCNRR:=5P8Hd>.RR;j2
F
OMN#0M80RHnP4dRUc:MRH0CCos=R:RC58b-0E442/ncdU;F
OMN#0M80RH4PUg:.RR0HMCsoCRR:=5b8C04E-24/Ug
.;O#FM00NMRP8HcnjgRH:RMo0CC:sR=8R5CEb0-/42cnjg;F
OMN#0M80RHjP.c:URR0HMCsoCRR:=5b8C04E-2j/.c
U;O#FM00NMRP8H4cj.RH:RMo0CC:sR=8R5CEb0-/424cj.;F
OMN#0M80RH4P6.RR:HCM0oRCs:5=R80CbE2-4/.64;O

F0M#NRM0LDFF6R4.:FRLFNDCM=R:RH58P.64Rj>R2O;
F0M#NRM0LDFF4cj.RL:RFCFDN:MR=8R5HjP4.>cRR;j2
MOF#M0N0FRLFjD.c:URRFLFDMCNRR:=5P8H.UjcRj>R2O;
F0M#NRM0LDFFcnjgRL:RFCFDN:MR=8R5HjPcg>nRR;j2
MOF#M0N0FRLF4DUg:.RRFLFDMCNRR:=5P8HU.4gRj>R2O;
F0M#NRM0LDFF4UndcRR:LDFFCRNM:5=R84HPncdURj>R2
;
O#FM00NMRl#k_8IH0:ERR0HMCsoCRR:=Apmm 'qhb5F#LDFF4+2RRmAmph q'#bF5FLFDR.2+mRAmqp hF'b#F5LF2DcRA+Rm mpqbh'FL#5FUFD2RR+Apmm 'qhb5F#LDFF4;n2
MOF#M0N0kR#lC_8bR0E:MRH0CCos=R:R-6RRm5Amqp hF'b#F5LF4D6.+2RRmAmph q'#bF5FLFD.4jc+2RRmAmph q'#bF5FLFDc.jU+2RRmAmph q'#bF5FLFDgcjn+2RRmAmph q'#bF5FLFDgU4.;22
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5kIl_HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_klI0H8E
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_b8C0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lC_8b20E;O

F0M#NRM0IH_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/OI_EOFHCH_I8R0E+;R4
MOF#M0N0_RI80CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E4I2/_FOEH_OC80CbERR+4
;
O#FM00NMRI8_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/8OHEFOIC_HE80R4+R;F
OMN#0M80R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/428E_OFCHO_b8C0+ERR
4;
MOF#M0N0_RI#CHxRH:RMo0CC:sR=_RII0H8Ek_MlC_ODRD#*_RI80CbEk_MlC_OD;D#
MOF#M0N0_R8#CHxRH:RMo0CC:sR=_R8I0H8Ek_MlC_ODRD#*_R880CbEk_MlC_OD;D#
F
OMN#0ML0RF_FD8RR:LDFFCRNM:5=R8H_#x-CRR#I_HRxC<j=R2O;
F0M#NRM0LDFF_:IRRFLFDMCNRR:=M5F0LDFF_;82
F
OMN#0MO0REOFHCH_I8R0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCH_I820E;F
OMN#0MO0REOFHCC_8bR0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCC_8b20E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8RI*5HE80-/428E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RRH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R5b8C04E-2_/8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IR5*R80CbE2-4/OI_EOFHCC_8b20ER4+R;-
-O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5855CEb0R4-R2RR/dR.2+5R55b8C0-ERRR42lRF8dR.2/nR42R2;R-R-RFyRVqR)vXd.4O1RC#DDRCMC8RC8
O--F0M#NRM0D0CV_CFPsRR:HCM0oRCs:5=R5C58bR0E+6R42FRl8.Rd2RR/4;n2RRRRRRRRRRRRRRRRRRRRRRRRRR--yVRFRv)q44nX1CRMC88CRsVFRVDC0PRFCIsRF#s8
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj4,RnH*I8_0EM_klODCD#6+4RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#nRR:F_k0L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNNDR8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDI8_N8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNNDR8osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2-;R-FR0RosCHC#0sER0CCR#D0CORo#HMRNDF0VRs0H#N
0CNs00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjjjj"RR&Ns8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjjjjj&"RR_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjRj"&8RN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
SRDRRFNI_8R8s<"=RjjjjjjjjjRj"&8RN_osC58dRF0IMF2Rj;C
SMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjj&"RR_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjj"jjRN&R8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjj"RR&Ns8_Cno5RI8FMR0Fj
2;S8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjj"RR&Ns8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj"jjRN&R8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjRj"&8RN_osC58gRF0IMF2Rj;C
SMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDI8_N8<sR=jR"j&"RR_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDI8_N8<sR=jR''RR&Ns8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R_N8s5Co48dRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;C
SMo8RCsMCNR0Cz;46
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzR4nRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0Rnz4;R
RR4Rz(:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2S;
CRM8oCCMsCN0R(z4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
pi-R-RR4Rzn:RRRRHV58N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HM-R-RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CM-R-RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;-R-RRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8bOsFC;##
S--CRM8oCCMsCN0Rnz4;-
-RRRRzR4(:VRHRF5M08RN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR_N8sRCo<q=R7;7)
S--CRM8oCCMsCN0R(z4;R
SR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1
4SzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>RcRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rc2<N=R8C_so85N8HsI8-0E4FR8IFM0R24c;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR4SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
-S-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.Sz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUX:4RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_ncdUX:4RRv)qA_4n1S4
RRRRRRRRRRRRb0FsRblNRQ575Rj2=H>RMC_so25[,7Rq7=)R>FRDI8_N84s5dFR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75Rj2=F>RkL0_k5#4H2,[2R;
RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRd<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;d2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRScz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..XRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gU4.RX.:qR)vnA4_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7R7)=D>RFNI_858s48.RF0IMF2Rj,hR RR=>',4'R)11RR=>',j'RS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm254RR=>F_k0L.k#5.H,*4[+27,Rm25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1Sc
zR.U:VRHRE5OFCHO_8IH0=ERRRc2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4R.2<N=R8C_so85N8HsI8-0E4FR8IFM0R24.;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzdRH:RVNR58I8sHE80R4>R.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;d4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgncRR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_cgcnXR):Rq4vAnc_1
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77RR=>D_FINs885R448MFI0jFR2 ,Rh>R=R''4,1R1)>R=R''j,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7dm52>R=R0Fk_#Lkc,5HR[c*+,d2R57m.=2R>kRF0k_L#Hc5,[c*+,.2RS
SSmS75R42=F>RkL0_k5#cH*,c[2+4,mR75Rj2=F>RkL0_k5#cHc,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5c[<2R=kRF0k_L#Hc5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*4[+2=R<R0Fk_#Lkc,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[.<2R=kRF0k_L#Hc5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+Rd2<F=RkL0_k5#cH*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d.
RRRRCRSMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_gz
Sd:dRRRHV5FOEH_OCI0H8ERR=go2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>4R42oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4R42<N=R8C_so85N8HsI8-0E4FR8IFM0R244;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUURR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_.cUUXR):Rq4vAng_1
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77RR=>D_FINs885R4j8MFI0jFR2 ,Rh>R=R''4,1R1)>R=R''j,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7(m52>R=R0Fk_#LkU,5HU+*[(R2,7nm52>R=R0Fk_#LkU,5HU+*[nR2,
SSSS57m6=2R>kRF0k_L#HU5,[U*+,62R57mc=2R>kRF0k_L#HU5,[U*+,c2R57md=2R>kRF0k_L#HU5,[U*+,d2RS
SSmS75R.2=F>RkL0_k5#UH*,U[2+.,mR75R42=F>RkL0_k5#UH*,U[2+4,mR75Rj2=F>RkL0_k5#UH*,U[R2,
SSSSu7Q5Rj2=H>RMC_so*5g[2+U,mR7u25jRR=>bHNs0L$_k5#UH2,[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5RH,[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>42jRRMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R24jRR<=Ns8_CNo58I8sHE80-84RF0IMFjR42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.XR4n:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv4cj.XR4n:qR)vnA4_U14
RSRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7R7)=D>RFNI_858sgFR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75246RR=>F_k0L4k#n,5H4[n*+246,mR7524cRR=>F_k0L4k#n,5H4[n*+24c,SR
S7SSmd542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm.542>R=R0Fk_#Lk4Hn5,*4n[.+427,Rm4542>R=R0Fk_#Lk4Hn5,*4n[4+42
,RSSSS74m5j=2R>kRF0k_L#54nHn,4*4[+jR2,7gm52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR75RU2=F>RkL0_kn#454H,n+*[U
2,SSSS7(m52>R=R0Fk_#Lk4Hn5,*4n[2+(,mR75Rn2=F>RkL0_kn#454H,n+*[nR2,76m52>R=R0Fk_#Lk4Hn5,*4n[2+6,S
SSRRRR57mc=2R>kRF0k_L#54nHn,4*c[+27,Rm25dRR=>F_k0L4k#n,5H4[n*+,d2R57m.=2R>kRF0k_L#54nHn,4*.[+2S,
SRRRRRRRR57m4=2R>kRF0k_L#54nHn,4*4[+27,Rm25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4u52>R=RsbNH_0$L4k#n,5HR[.*+,42Ru7m5Rj2=b>RN0sH$k_L#54nH.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_dSn
zRcd:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>RRg2CRoMNCs0SC
RRRRz	OD:sRbF#OC#BR5p
i2SRSRLHCoMS
SRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSSRRRRRsN8CNo58I8sHE80-84RF0IMF2RgRR<=Ns8_CNo58I8sHE80-84RF0IMF2Rg;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RSRRcRzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSz6RR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SSsSI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0Cz;c6
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SSnzcRH:RVNR58I8sHE80RR<=go2RCsMCN
0CSSSSF_k0CHM52=R<R''4;S
SSsSI0M_C5RH2<W=R S;
SMSC8CRoMNCs0zCRc
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#S
SS(zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.d:.RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRARR)_qv6X4.d:.RRv)qA_4n1
dnRRRRRRRRRRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cdo5n+*[d84RF0IMFnRd*,[2R7q7)>R=D_FINs8858URF0IMF2Rj,hR RR=>',4'R)11RR=>',j'
RRRRRRRRRRRRRRRRRRRRRRRRRRRRWRR >R=R0Is_5CMHR2,BRpi=B>RpRi,7dm54=2R>kRF0k_L#5d.H.,d*d[+4R2,7dm5j=2R>kRF0k_L#5d.H.,d*d[+j
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR752.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR752.(RR=>F_k0Ldk#.,5Hd[.*+2.(,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5n=2R>kRF0k_L#5d.H.,d*.[+nR2,7.m56=2R>kRF0k_L#5d.H.,d*.[+6R2,7.m5c=2R>kRF0k_L#5d.H.,d*.[+c
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR752..RR=>F_k0Ldk#.,5Hd[.*+2..,mR752.4RR=>F_k0Ldk#.,5Hd[.*+2.4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5j=2R>kRF0k_L#5d.H.,d*.[+jR2,74m5g=2R>kRF0k_L#5d.H.,d*4[+gR2,74m5U=2R>kRF0k_L#5d.H.,d*4[+U
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR75246RR=>F_k0Ldk#.,5Hd[.*+246,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR74m5c=2R>kRF0k_L#5d.H.,d*4[+cR2,74m5d=2R>kRF0k_L#5d.H.,d*4[+dR2,74m5.=2R>kRF0k_L#5d.H.,d*4[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4542>R=R0Fk_#LkdH.5,*d.[4+427,Rmj542>R=R0Fk_#LkdH.5,*d.[j+427,Rm25gRR=>F_k0Ldk#.,5Hd[.*+,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Um52>R=R0Fk_#LkdH.5,*d.[2+U,mR75R(2=F>RkL0_k.#d5dH,.+*[(R2,7nm52>R=R0Fk_#LkdH.5,*d.[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m6=2R>kRF0k_L#5d.H.,d*6[+27,Rm25cRR=>F_k0Ldk#.,5Hd[.*+,c2R57md=2R>kRF0k_L#5d.H.,d*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75R.2=F>RkL0_k.#d5dH,.+*[.R2,74m52>R=R0Fk_#LkdH.5,*d.[2+4,mR75Rj2=F>RkL0_k.#d5dH,.2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,75mud=2R>NRbs$H0_#LkdH.5,*Rc[2+d,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mu.=2R>NRbs$H0_#LkdH.5,*Rc[2+.,mR7u254RR=>bHNs0L$_k.#d5RH,c+*[4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u25jRR=>bHNs0L$_k.#d5RH,c2*[2R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSCRM8oCCMsCN0R(zc;S
SCRM8oCCMsCN0Rczc;C
SMo8RCsMCNR0Cz;cd
8CMRONsECH0Os0kCFRM__sIOOEC	
;
---
-NRp#H0RlCbDl0CMNF0HM#RHRV8CN0kD

--NEsOHO0C0CksRD#CC_O0sRNlF)VRq)v_WHuR#k
VMHO0FoMRCC0_M88_CEb05x#HCRR:HCM0oRCs;CR8bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCHRlMH_#x:CRR0HMCsoCRR:=jL;
CMoH
lRRH#M_HRxC:8=RCEb0;R
RH5VR#CHxR8<RCEb02ER0CRM
RlRRH#M_HRxC:#=RH;xC
CRRMH8RVR;
R0sCkRsMl_HM#CHx;M
C8CRo0M_C8C_8b;0E
MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R855CEb0R4-R2n/42R;RRRRRRRRRR-R-RFyRVqR)vX4n4O7RC#DDRCMC8
C80C$bR0Fk_#Lk_b0$C#RHRsNsN5$RM_klODCD#FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k:#RR0Fk_#Lk_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COFds5RI8FMR0FjR2;RRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD8RN8#s_0:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--bCHbDCHMRNsC8CRso0H#CNs
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80Rc<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRR4:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&8RN8#s_0jo52R;
RRRRRDRRFII_Ns88RR<="jjj"RR&Ns8_Cjo52R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=RjRj"&8RN8#s_04o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&Ns8_C4o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&8RN8#s_0.o5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R''jRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E>2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<N=R8_8s#50odFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=8RN_osC58dRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRc
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR6:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR6R;
RzRRn:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rh7Q;R
RRMRC8CRoMNCs0zCRn
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR(RzRRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soL2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC;R
RRMRC8CRoMNCs0zCRU
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
R--RzRRg:RRRRHV58N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HM-R-RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CM-R-RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;-R-RRRRRRRRRRMRC8VRH;-
-RRRRRRRRCRM8bOsFC;##
R--RCRRMo8RCsMCNR0Cz
g;-R-RR4RzjRR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)-;
-RRRR8CMRMoCC0sNC4RzjR;
RRRRR
RRRRRR-b-RHDbCHRMC#o0NCs8RC#oH0
CsRRRRzR46Rb:RsCFO#5#RB,piR_N8s2Co
RSRRoLCHRM
RRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRR8N8s0_#o=R<R_N8s5CoNs88I0H8ER-48MFI0jFR2R;
RRRRRCRRMH8RVR;
RCRRMb8RsCFO#z#R4
6;RRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR44:FRVsRRHHMMRkOl_C#DDRI8FMR0FjCRoMNCs0RC
RRRRR-RR-VRQR85N8HsI8R0E>2RcRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4.:VRHR85N8HsI8R0E>2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58N8s0_#o85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI0cFR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rz.R;
RRRRR-RR-VRQR85N8HsI8R0E<c=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:dRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC4RzdR;
R-RR-MRtC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:cRRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)Rqv:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4Rn2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR):qvRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds527,Ruj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42RR
RRRRRRRRRRRRRRRRRRRRRRRRR7qu).>R=RIDF_8sN8.s527,Rud)qRR=>D_FIs8N8s25d, RWRR=>I_s0CHM52
,RRRRRRRRRRRRRRRRRRRRRRRRRRBRWp=iR>pRBi7,Ru=mR>kRF0k_L#,5H[;22
RRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_kH#5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR
MN8RsHOE00COkRsC#CCDOs0_N
l;
