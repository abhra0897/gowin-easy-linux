--
@ER--RbBF$osHE50RO42RgRgg1b$MDHHO0R$,Q3MO
R--RDqDRosHER0#sCC#s8PC3-
-
R--#CCDOF0HMCR#0CR8VHHM0MHF3WRRCHRIDCDRP0CMkDND$8RN8DRLF_O	sRFl0
FF-N-RsDOEHR#0=CR#D0CO_lsF

---f-R]8CNCRs:/$/#MHbDO$H0/blN.N4.OlG/NCbbsG#/HMDHGH/DLC/oMb_#NNs0Msd/FPl3E48yR-f
-D

HNLssH$RC;CC
#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCFRIso	3CNMbOo	NCD3ND
;
DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$)_mvLCN#R
H#SMoCCOsHRS5
SHSI8R0E:MRH0CCos=R:R
c;SNSS8I8sHE80RH:RMo0CC:sR=;R(
SSSDNFI8R8s:MRH0CCos=R:R
j;SESSHNoE8R8s:MRH0CCos=R:R;(U
SSS0DNLCRR:s0FlNCLD;S
SSD8V0RR:sIFlF
s8S
2;SsbF0
R5SqSS7R7):MRHR8#0_oDFHPO_CFO0sNR58I8sHE80R4-RRI8FMR0Fj
2;S7SSmRza:kRF00R#8F_Do_HOP0COF5sRI0H8ERR-4FR8IFM0R
j2S;S2
0SN0LsHkR0CQahQR#:R0MsHoS;
Ns00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;CRM8CHM00)$RmLv_N;#C
s
NO0EHCkO0s#CRCODC0m_)vVRFRv)m_#LNC#RH
kS#Lb0$CFRsl0FkRRH##_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;-O-SFFlbM0CMRXvzw-n
-bSSFRs05-
-SSSSm:RRR0FkR8#0_oDFH
O;-S-SSjSQRH:RM0R#8F_Do;HO
S--SQSS4RR:H#MR0D8_FOoH;-
-SSSS1:RRRRHM#_08DHFoO-
-S2SS;-
-S8CMRlOFbCFMMS0;
O
SF0M#NRM0ERCG:0R#soHM50jRF6R42=R:R4"j.6dcng(Uq7AB ;w"
V
Sk0MOHRFMs0FlNCLDs8CN5L0ND:CRRlsF0DNLCI;R,,RLRMDCRH:RMo0CCRs2skC0s#MR0MsHo>R=RF"slL0NDCCsN;8"
V
Sk0MOHRFMVOkMP5NDL0F0FHlDMVC_,FRDI8N8s,_VRoEHE8N8s,_VR0LH,LRMHR0#:MRH0CCoss2RCs0kM0R#soHMR
H#SFSOMN#0M00RF:bRR0HMCsoCRR:=L0F0FHlDMVC_RM+RL#H0R4-R;S
SPHNsNCLDRRH,[P,R,bRLF:#RR0HMCsoC;S
SO#FM00NMRb0FOsENRH:RMo0CC:sR=LRMHR0#/RRc-;R4
PSSNNsHLRDCLRkV:0R#soHM5b0FOsENRI8FMR0Fj
2;SoLCHSM
S5HVL0F0FHlDMVC_RD<RF8IN8Vs_RRFs0RFb>HREo8EN8Vs_2ER0CSM
SRS[:j=R;S
SS:PR=;Rj
SSSL#bFRR:=jS;
SFSVsRRHHLMRFF00lMDHCR_V00FRFRbRDbFF
SSSSRHVHRR<DNFI8_8sVsRFR>HRRoEHE8N8sR_V0MEC
SSSSVSHRD8V0H5L0=2RR''4RC0EMS
SSSSSP=R:R+PRR*.*[S;
SSSSCRM8H
V;SSSSCCD#
SSSSVSHRL0NDHC52H5L0=2RR''4RC0EMS
SSSSSP=R:R+PRR*.*[S;
SSSSCRM8H
V;SSSSCRM8H
V;SSSS[=R:R+[RRR4;R-RR-kRMlsLCRRFVL#H0RDOFD0COC
8RSSSSH[V5Rc=R2ER0C-MR-PRCCRs$cCRIRl8kbMRH0NFRRNOEs0NOCSs
SSSS[=R:R
j;SSSSSVLk5FLb#:2R=CREG25P;S
SSLSSbRF#:L=RbRF#+;R4
SSSSRSP:j=R;S
SSMSC8VRH;S
SS8CMRFDFbS;
SCSs0MksRVLk;S
SCCD#
SSSskC0ssMRFNl0LsDCC5N80DNLCL,RFF00lMDHC,_VR0LH,LRMH20#;S
SCRM8H
V;S8CMRMVkOF0HMkRVMNOPD
;
SMOF#M0N0FRL0l0FpCHMRH:RMo0CC:sR=DR5F8IN84s/n42*nS;
O#FM00NMR0LF0dFl.MpHCRR:HCM0oRCs:5=RDNFI8/8sd*.2d
.;SMOF#M0N0HREoHEpM:CRR0HMCsoCRR:=5oEHE8N8sn/42n*4;O
SF0M#NRM0EEHodH.pM:CRR0HMCsoCRR:=5oEHE8N8s./d2.*d;O
SF0M#NRM0EEHoA8FsC:sRR0HMCsoCRR:=EEHopCHMR4+R6
R;SMOF#M0N0sR0HN#00HC_RH:RMo0CC:sR=ER5HAoEFCs8s-+4L0F0FHlpM/C24;nR
$S0b0CRNHLR#sRNsRN$5H5Eo.EdpCHMRL-RFF00lpd.H2MC/+d.4FR8IFM0RRj2FsVRFklF0
R;So#HMRND1amz,mRpz:aRRL0N;#
SHNoMDmR7zNa_kRG,7amz_GNk.RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;LHCoMR
RRVRRFbs_H:bCRsVFRHHRMRRj0IFRHE80-o4RCsMCN
0CS0SN0LsHkR0C\N3sMR	\FsVRCRo#:NRDLRCDH4#R;R
RRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;SCRLo
HMSsSRC:o#RbbHCVLk
SSSRsbF0NRlbS5
RSRRSRSSR=QR>mR7zNa_kHG52S,
RSRRSRSSR=mR>mR7zHa52S
SSRSS2S;
R8CMRMoCC0sNCFRVsH_bb
C;
VSH_#4n:VRHRH5Eo.EdpCHMRL>RFF00lpd.H2MCRMoCC0sNCS
SLHCoMS
SH4V_nRL:H5VRL0F0FHlpM=CRR0LF0dFl.MpHCo2RCsMCN
0CSLSS:FRVsHRL0MRHR0jRFHRI8R0E-RR4oCCMsCN0
SSSS0N0skHL0QCRhRQaF)VRm6v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,d;.2
SSSLHCoMS
SSmS)vR 6:mR)vXd.4S
SSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSq=cR>7Rq7c)52S,
SSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SMSC8CRoMNCs0LCR;S
SCRM8oCCMsCN0R_HV4;nL
HSSVn_4LH:RVLR5FF00lMpHCRR>L0F0F.ldpCHM2CRoMNCs0SC
S:SLRsVFR0LHRRHMjFR0R8IH0-ERRo4RCsMCN
0CSSSSNs00H0LkChRQQFaRVmR)vR c:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SLSSCMoH
SSSSv)m :cRRv)m44nX
SSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSqSS4>R=R7q7)254,S
SSSSSSqSS.>R=R7q7)25.,S
SSSSSSqSSd>R=R7q7)25d,S
SSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SS8CMRMoCC0sNC;RL
CSSMo8RCsMCNR0CH4V_n
L;S8CMRMoCC0sNCVRH_#4n;S

HdV_.R#:H5VREEHodH.pM=CRR0LF0dFl.MpHCo2RCsMCN
0CSVSH_O4n:VRHRF5L0l0FpCHMRL=RFF00lpd.H2MCRMoCC0sNCS
SSRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SHSSV:_4RRHV58N8s8IH0=ERRR42oCCMsCN0
SSSS0SN0LsHkR0CQahQRRFV) mv4RR:DCNLD#RHRMVkODPN50LF0pFlH,MCRIDFNs88,HREo8EN8Rs,L,H0R24n;S
SSCSLo
HMSSSSSv)m :4RRv)m44nX
SSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSSRq4='>Rj
',SSSSSSSSS.SqRR=>',j'
SSSSSSSSqSSd>R=R''j,S
SSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSS2S;
SCSSMo8RCsMCNR0CH4V_;S
SSVSH_R.:H5VRNs88I0H8ERR=.o2RCsMCN
0CSSSSS0N0skHL0QCRhRQaF)VRm.v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSoLCHSM
SSSS) mv.RR:)4mvn
X4SSSSSbSSFRs0lRNb5qRRj>R=R7q7)25j,S
SSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSSRq.='>Rj
',SSSSSSSSSdSqRR=>',j'
SSSSSSSSmSSR>R=Rz1ma25j50LH2S
SSSSSS2SS;S
SSMSC8CRoMNCs0HCRV;_.
SSSS_HVdH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
SSSSNs00H0LkChRQQFaRVmR)vR d:NRDLRCDHV#RkPMONLD5FF00lMpHCD,RF8IN8Rs,EEHoNs88,HRL04,Rn
2;SSSSLHCoMS
SS)SSmdv R):Rmnv4XS4
SSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSRqd='>Rj
',SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSS2S;
SCSSMo8RCsMCNR0CHdV_;S
SSVSH_Rc:H5VR5oEHE8N8sF-L0l0FpCHMR4<RnN2RM58RNs88I0H8E=R>R2c2RMoCC0sNCS
SSNSS0H0sLCk0RQQhaVRFRv)m :cRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SLSSCMoH
SSSSmS)vR c:mR)vX4n4S
SSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSSRmR=1>Rm5zajL25H
02SSSSSSSSS
2;SSSSCRM8oCCMsCN0R_HVcS;
SHSSV:_6RRHV585N8HsI8R0E>6=R2MRN8ER5HNoE8R8s-FRL0l0FpCHMRR>=42n2RMoCC0sNCS
SSNSS0H0sLCk0RQQhaVRFRv)m :6RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,.Rd2S;
SLSSCMoH
SSSSmS)vR 6:mR)vXd.4S
SSSSSSsbF0NRlbRR5RRqj=q>R757)j
2,SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSqSS.>R=R7q7)25.,S
SSSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSSRqc=q>R757)c
2,SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS;S2
SSSS8CMRMoCC0sNCVRH_
6;SCSSMo8RCsMCNR0CLS;
S8CMRMoCC0sNCVRH_O4n;S
SH4V_nR8:H5VRL0F0FHlpM>CRR0LF0dFl.MpHCo2RCsMCN
0CSHSSV8_Ns8IH0RE:H5VRNs88I0H8ERR>co2RCsMCN
0CSSSSLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SSHSSV:_cRRHV5H5Eo8EN8Ls-FF00lMDHCRR<4Rn2NRM858N8s8IH0>ER=2Rc2CRoMNCs0SC
SSSSS0N0skHL0QCRhRQaF)VRmcv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSCSLo
HMSSSSSmS)vR c:mR)vX4n4S
SSSSSSFSbsl0RN5bRRRqj=q>R757)j
2,SSSSSSSSSqSS4>R=R7q7)254,S
SSSSSSSSSSRq.=q>R757).
2,SSSSSSSSSqSSd>R=R7q7)25d,S
SSSSSSSSSS=mR>mR1zja52H5L0S2
SSSSSSSSS;S2
SSSSMSC8CRoMNCs0HCRV;_c
SSSS8CMRMoCC0sNC;RL
SSSCRM8oCCMsCN0R_HVNI8sHE80;S
SS_HVNs88I0H8EH:RVNR58I8sHE80RR<=co2RCsMCN
0CSSSSLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SSHSSV:_4RRHV58N8s8IH0=ERRR42oCCMsCN0
SSSSNSS0H0sLCk0RQQhaVRFRv)m :4RRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SSSSLHCoMS
SSSSS) mv4RR:)4mvn
X4SSSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSS4SqRR=>',j'
SSSSSSSSSSSq=.R>jR''S,
SSSSSSSSSdSqRR=>',j'
SSSSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSSSSSS
2;SSSSS8CMRMoCC0sNCVRH_
4;SSSSS_HV.H:RVNR58I8sHE80R.=R2CRoMNCs0SC
SSSSS0N0skHL0QCRhRQaF)VRm.v RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSCSLo
HMSSSSSmS)vR .:mR)vX4n4S
SSSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSS.SqRR=>',j'
SSSSSSSSSSSq=dR>jR''S,
SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS2SS;S
SSCSSMo8RCsMCNR0CH.V_;S
SSHSSV:_dRRHV58N8s8IH0=ERRRd2oCCMsCN0
SSSSNSS0H0sLCk0RQQhaVRFRv)m :dRRLDNCHDR#kRVMNOPDF5L0l0FpCHM,FRDI8N8sE,RHNoE8,8sR0LH,nR42S;
SSSSLHCoMS
SSSSS) mvdRR:)4mvn
X4SSSSSSSSb0FsRblNRR5Rq=jR>7Rq7j)52S,
SSSSSSSSS4SqRR=>q)775,42
SSSSSSSSSSSq=.R>7Rq7.)52S,
SSSSSSSSSdSqRR=>',j'
SSSSSSSSSSSm=RR>mR1zja52H5L0S2
SSSSS2SS;S
SSCSSMo8RCsMCNR0CHdV_;S
SSHSSV:_cRRHV5H5Eo8EN8Ls-FF00lMDHCRR<4Rn2NRM858N8s8IH0>ER=2Rc2CRoMNCs0SC
SSSSS0N0skHL0QCRhRQaF)VRmcv RD:RNDLCRRH#VOkMP5NDL0F0FHlpMRC,DNFI8,8sRoEHE8N8sL,RHR0,4;n2
SSSSCSLo
HMSSSSSmS)vR c:mR)vX4n4S
SSSSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSSSSq=4R>7Rq74)52S,
SSSSSSSSS.SqRR=>q)775,.2
SSSSSSSSSSSq=dR>7Rq7d)52S,
SSSSSSSSSRSmRR=>1amz55j2L2H0
SSSSSSSS
2;SSSSS8CMRMoCC0sNCVRH_
c;SSSSCRM8oCCMsCN0R
L;SCSSMo8RCsMCNR0CHNV_8I8sHE80;S
SCRM8oCCMsCN0R_HV4;n8
MSC8CRoMNCs0HCRV._d#
;
S:L4RsVFRHIRMRR405FREEHodH.pM-CRR0LF0dFl.MpHC.-d2./dRMoCC0sNCS
SLV:RFLsRHH0RMRRj0IFRHE80R4-RRMoCC0sNCS
SS0N0skHL0QCRhRQaF)VRm6v RD:RNDLCRRH#VOkMP5NDI.*d+0LF0dFl.MpHCD,RF8IN8Rs,EEHoNs88,HRL0d,R.
2;S#SSHNoMDHRbb8C_F#k0R#:R0D8_FOoH;S
SLHCoMS
SSv)m :6RRv)md4.X
SSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSRq4=q>R757)4
2,SSSSSSSSq=.R>7Rq7.)52S,
SSSSSqSSd>R=R7q7)25d,S
SSSSSScSqRR=>q)775,c2
SSSSSSSSRmR=1>Rm5zaIL25H
02SSSSS2SS;S
SCRM8oCCMsCN0R
L;S8CMRMoCC0sNC4RL;S

H4V_nRF:H5VR5oEHEpd.HRMC=ERRHpoEH2MCR8NMRH5Eo.EdpCHMRL>RFF00lpd.H2MC2CRoMNCs0SC
SRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SHS#oDMNR0Fk_8CMR#:R0D8_FOoH;S
SS0N0skHL0QCRhRQaF)VRmcv RD:RNDLCRRH#VOkMP5NDEEHoA8FsC4s-6E,RHAoEFCs8s6-4,HREo8EN8Rs,L,H0R24n;S
SLHCoMS
SSv)m :cRRv)m44nX
SSSSFSbsl0RN5bRRRqjRR=>q)775,j2
SSSSSSSSRq4=q>R757)4
2,SSSSSSSSq=.R>7Rq7.)52S,
SSSSSqSSd>R=R7q7)25d,S
SSSSSSRSmRR=>1amz5H5Eo.EdpCHM-0LF0dFl.MpHC.-d2./d+542L2H0
SSSSSSS2S;
S8CMRMoCC0sNC;RL
MSC8CRoMNCs0HCRVn_4FS;
H4V_nR#:H5VR5oEHEpd.HRMC<ERRHpoEH2MCR8NMRH5Eo.EdpCHMRL>RFF00lpd.H2MC2CRoMNCs0SC
SRL:VRFsLRH0HjMRRR0FI0H8ERR-4CRoMNCs0SC
SHS#oDMNR0Fk_8CMR#:R0D8_FOoH;S
SS0N0skHL0QCRhRQaF)VRm6v RD:RNDLCRRH#VOkMP5NDEEHoA8FsCds-4E,RHAoEFCs8s4-d,HREo8EN8Rs,L,H0R2d.;S
SLHCoMS
SSv)m :6RRv)md4.X
SSSSFSbsl0RN5bRRjRqRR=>q)775,j2
SSSSSSSSRq4=q>R757)4
2,SSSSSSSSq=.R>7Rq7.)52S,
SSSSSqSSd>R=R7q7)25d,S
SSSSSScSqRR=>q)775,c2
SSSSSSSSRmR=1>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM2./d2H5L0S2
SSSSS;S2
CSSMo8RCsMCNR0CLS;
CRM8oCCMsCN0R_HV4;n#
R
RRVRH_8IH0RE:H5VR0#sH0CN0_<HRRR62oCCMsCN0
RRRRRRRR_HVFjk0:VRHRH5Eo.EdpCHMRL=RFF00lpd.H2MCRMoCC0sNCR
RRRRRRRRRRzpma25jRR<=1amz5;j2
RRRRRRRR8CMRMoCC0sNCVRH_0FkjR;
RRRRRHRRVk_F0R4:H5VREEHodH.pM>CRR0LF0dFl.MpHCo2RCsMCN
0CRRRRRRRRRHRRVN_O#:C4RRHV50LF0pFlHRMC=FRL0l0FdH.pMRC2oCCMsCN0
S--So#HMRND8VHVR#:R0D8_FOoH;R
SRCRLo
HM-R-RRRRRRRRRRRRR8VHVRR<='Rj'IMECR7q7)=R<RhBmea_17m_pt_QBea Bmd)54F+L0l0FpCHM,8RN8HsI820ER-
-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDC4R''-;
-RSRRRRRV_FsI0H8EV:RFHsRRRHMjFR0R8IH04E-RMoCC0sNC-
-SRRRRRRRRkRlGC0sCRR:vwzXn-
-SbSSFRs0lRNb5-
-SSSSRRRmRR=>pamz55j2H
2,-S-SSRSRQ=jR>mR1zja5225H,-
-SSSSR4RQRR=>1amz5542H
2,-S-SSRSR1=RR>HR8V-V
-SSS2-;
-RRRRRRRRRRRRCRRMo8RCsMCNR0CV_FsI0H8ER;
RRRRRRRRRRRRRzpma25jRR<=1amz5Rj2IMECR7q7)=R<RhBmea_17m_pt_QBea Bmd)54F+L0l0FpCHM,8RN8HsI820ERR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C1amz5;42
RRRRRRRRRRRCRM8oCCMsCN0R_HVOCN#4R;
RRRRRRRRRVRH_#ONCR.:H5VRL0F0FHlpM>CRR0LF0dFl.MpHCo2RCsMCN
0C-S-S#MHoN8DRHjVVR#:R0D8_FOoH;R
SRLRRCMoH
R--RRRRRRRRRRRRRV8HV<jR=jR''ERICqMR7R7)<B=Rm_he1_a7pQmtB _eB)am5+46L0F0FHlpMRC,Ns88I0H8E
2R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#'CR4
';-R-SRRRRRsVF_8IH0:EjRsVFRHHRMRRj0IFRHE80-o4RCsMCN
0C-R-SRRRRRRRRl0kGsRCC:zRvX
wn-S-SSsbF0NRlb
R5-S-SSRSRm=RR>mRpzja5225H,-
-SSSSRjRQRR=>1amz55j2H
2,-S-SSRSRQ=4R>mR1z4a5225H,-
-SSSSRRR1RR=>8VHVj-
-S2SS;-
-RRRRRRRRRRRRRMRC8CRoMNCs0VCRFIs_HE80jR;
RRRRRRRRRRRRRzpma25jRR<=1amz5Rj2IMECR7q7)=R<RhBmea_17m_pt_QBea Bm4)56F+L0l0FpCHM,8RN8HsI820ERR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C1amz5;42
RRRRRRRRRRRCRM8oCCMsCN0R_HVOCN#.R;
RRRRRCRRMo8RCsMCNR0CHFV_k;04
RRRRRRRRRN:VRFsIMRHR04RFER5HdoE.MpHCRR-L0F0F.ldpCHM-2d./-d.4CRoMNCs0-C
-#SSHNoMDHR8VRV4:0R#8F_Do_HOP0COF5s5EEHodH.pM-CRR0LF0dFl.MpHC.-d2./d-84RF0IMF2R4;R
SRLRRCMoH
R--RRRRRRRRRRRRRV8HVI452=R<R''jRCIEM7Rq7<)RRhBmea_17m_pt_QBea Bmd)5.I*5++42L0F0F.ldpCHM,8RN8HsI820E
R--RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#R''4;-
-SRRRRVRRFIs_HE804V:RFHsRRRHMjFR0R8IH04E-RMoCC0sNC-
-SRRRRRRRRkRlGC0sCRR:vwzXn-
-SbSSFRs0lRNb5-
-SSSSRRRmRR=>pamz55I2H
2,-S-SSRSRQ=jR>mRpzIa5-542H
2,-S-SSRSRQ=4R>mR1zIa5+542H
2,-S-SSRSR1=RR>HR8V5V4I-2
-SSS2-;
-RRRRRRRRRRRRCRRMo8RCsMCNR0CV_FsI0H8E
4;RRRRRRRRRRRRRmRpzIa52=R<Rzpma-5I4I2RERCMq)77RB<Rm_he1_a7pQmtB _eB)am5*d.54I+2F+L0l0FdH.pMRC,Ns88I0H8ER2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#Rz1ma+5I4
2;RRRRRRRRCRM8oCCMsCN0R
N;RRRRRRR
RRRRRHRRVN_D#n04:VRHRE55HdoE.MpHCRR=EEHopCHM2MRN8ER5HdoE.MpHCRR-L0F0F.ldpCHMRn>RdR22oCCMsCN0
S--So#HMRND8VHV.RR:#_08DHFoOS;
RRRRLHCoM-
-RRRRRRRRRRRRRHR8VRV.<'=RjI'RERCMq)77RB<Rm_he1_a7pQmtB _eB)am5oEHEsAF8-Cs4R6,Ns88I0H8E
2R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C';4'
S--RRRRRFRVsH_I8.0E:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
S--RRRRRRRRRGlk0CsCRv:RznXw
S--SFSbsl0RN5bR
S--SRSSRRmR=p>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./2d.5,H2
S--SRSSRRQj=p>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./-d.4H252-,
-SSSSQRR4>R=Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2d5.2H
2,-S-SSRSR1=RR>HR8V
V.-S-SS
2;-R-RRRRRRRRRRRRRCRM8oCCMsCN0RsVF_8IH0;E.
RRRRRRRRRRRRzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.<2R=mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d4.-2SR
SSSSIMECR7q7)RR<Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,46R8N8s8IH0
E2RRRRRRRRRRRRRRRRRRRRCCD#Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2d;.2
RRRRRRRR8CMRMoCC0sNCVRH_#DN0;4n
R
RRRRRRVRH_#DN0:d.RRHV5H5Eo.EdpCHMRR<REEHopCHM2MRN8ER5HdoE.MpHCRR-L0F0F.ldpCHMRn>RdR22oCCMsCN0
S--So#HMRND8VHVdRR:#_08DHFoOS;
RRRRLHCoM-
-RRRRRRRRRRRRRHR8VRVd<'=RjI'RERCMq)77RB<Rm_he1_a7pQmtB _eB)am5oEHEsAF8-CsdR4,Ns88I0H8E
2R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#C';4'
S--RRRRRFRVsH_I8d0E:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
S--RRRRRRRRRGlk0CsCRv:RznXw
S--SFSbsl0RN5bR
S--SRSSRRmR=p>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./2d.5,H2
S--SRSSRRQj=p>Rm5za5oEHEpd.H-MCL0F0F.ldpCHM-2d./-d.4H252-,
-SSSSQRR4>R=Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2d5.2H
2,-S-SSRSR1=RR>HR8V
Vd-S-SS
2;-R-RRRRRRRRRRRRRCRM8oCCMsCN0RsVF_8IH0;Ed
RRRRRRRRRRRRzpmaE55HdoE.MpHCF-L0l0FdH.pMdC-.d2/.<2R=mRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d4.-2SR
SSSSIMECR7q7)RR<Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C-,d4R8N8s8IH0
E2RRRRRRRRRRRRRRRRRRRRCCD#Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2d;.2
RRRRRRRR8CMRMoCC0sNCVRH_#DN0;d.
R
RRRRRRVRH_0Fk.H:RVER5HAoEFCs8sRR-L0F0FHlpM<CRR2ncRMoCC0sNCR
RRRRRRRRRRRRR7amz_GNkRR<=80VDRCIEMRR5R5RRq)77RB>Rm_he1_a7pQmtB _eB)am5oEHEsAF8,CsR8N8s8IH02E2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRFR75q7<)RRhBmea_17m_pt_QBea BmL)5FF00lMpHCN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#Cpamz5;j2
RRRRRRRR8CMRMoCC0sNCVRH_0Fk.R;
RRRRRHRRVk_F0Rd:H5VREEHoA8FsC-sRR0LF0pFlHRMC>dRn2CRoMNCs0RC
RRRRRRRRRRRRRz7mak_NG=R<RD8V0ERIC5MRRRRR57q7)RR>Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRF5sRq)77RB<Rm_he1_a7pQmtB _eB)am50LF0pFlH,MCR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRR#CDCmRpz5a5EEHodH.pMLC-FF00lpd.H-MCd/.2d;.2
RRRRRRRR8CMRMoCC0sNCVRH_0FkdR;
RRRRCRM8oCCMsCN0R_HVI0H8ER;
RRR
RRRRHIV_HE80jH:RV0R5s0H#N_0CH=R>RR62oCCMsCN0
RRRRRRRR_HVOCN#4H:RVLR5FF00lMpHCRR=L0F0F.ldpCHM2CRoMNCs0RC
RRRRRRRRRmR7zNa_k<GR=mR1zja52ERIC5MRRRRR57q7)=R<RhBmea_17m_pt_QBea Bmd)54F+L0l0FpCHM,8RN8HsI820E2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRM857q7)=R>RhBmea_17m_pt_QBea BmL)5FF00lMpHCN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HVOCN#4R;
RRRRRHRRVN_O#:C.RRHV50LF0pFlHRMC>FRL0l0FdH.pMRC2oCCMsCN0
RRRRRRRRRRR7amz_GNkRR<=1amz5Rj2IMECRR5RRqR57R7)<B=Rm_he1_a7pQmtB _eB)am5+46L0F0FHlpMRC,Ns88I0H8ER22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSNRM857q7)=R>RhBmea_17m_pt_QBea BmL)5FF00lMpHCN,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HVOCN#.R;
RRRRRNRRjV:RFIsRRRHM4FR0RH5Eo.EdpCHM-0LF0dFl.MpHC.-d2./dRMoCC0sNCR
RRRRRRRRRRRRR7amz_GNkRR<=1amz5RI2IMECRR5RRqR57R7)<B=Rm_he1_a7pQmtB _eB)am5*d.54I+2L+RFF00lpd.H-MC4N,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRRM58Rq)77RR>=Bemh_71a_tpmQeB_ mBa).5d*LI+FF00lpd.H,MCR8N8s8IH02E22R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCjRN;R
RRRRRRVRH_b#kdR.:H5VR5oEHEpd.HRMC=ERRHpoEH2MCR8NMRH5Eo.EdpCHMRL-RFF00lpd.HRMC>dRn2o2RCsMCN
0CRRRRRRRRRRRRRmR7zNa_k<GR=mR1z5a5EEHodH.pMLC-FF00lpd.H2MC/2d.RS
SSSRRSISSERCM5RRRR75q7<)R=mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCRs,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRN8qR57R7)>B=Rm_he1_a7pQmtB _eB)am5oEHEsAF8-Cs4R6,Ns88I0H8E222
RRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCFRsl0Fk'05FE#CsRR=>'2Z';R
RRRRRRMRC8CRoMNCs0HCRVk_#b;d.
RRRRRRRR_HV#4kbnH:RV5R5EEHodH.pM<CRRHREoHEpMRC2NRM85oEHEpd.HRMC-FRL0l0FdH.pM>CRR2nd2CRoMNCs0RC
RRRRRRRRRRRRRz7mak_NG=R<Rz1maE55HdoE.MpHCF-L0l0FdH.pM/C2dR.2
SSSRSRSSESIC5MRRRRR57q7)=R<RhBmea_17m_pt_QBea BmE)5HAoEFCs8sN,R8I8sHE802R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8NMR75q7>)R=mRBh1e_ap7_mBtQ_Be a5m)EEHoA8FsCds-4N,R8I8sHE802
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RlsFF'k05EF0CRs#='>RZ;'2
RRRRRRRR8CMRMoCC0sNCVRH_b#k4
n;RRRRRRRRHDV_FRI:H5VRL0F0FHlpM>CRRRj2oCCMsCN0
RRRRRRRRRRR7amz_GNkRR<=80VDRCIEMRR5RqR57R7)<mRBh1e_ap7_mBtQ_Be a5m)L0F0FHlpMRC,Ns88I0H8E
22RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRSRRFs57q7)RR>Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R2
RRRRRRRRRRRRRRRRRRRRRCRRDR#CsFFlk50'FC0Es=#R>ZR''
2;RRRRRRRRCRM8oCCMsCN0R_HVD;FI
RRRRRRRR_HVDjFI:VRHRF5L0l0FpCHMR4<R2CRoMNCs0RC
RRRRRRRRRmR7zNa_k<GR=VR8DI0RERCM57q7)RR>Bemh_71a_tpmQeB_ mBa)H5EoFEAss8C,8RN8HsI820E2R
RRRRRRRRRRRRRRRRRRRRRRDRC#sCRFklF0F'50sEC#>R=R''Z2R;
RRRRRCRRMo8RCsMCNR0CHDV_F;Ij
RRRRMRC8CRoMNCs0HCRVH_I8j0E;C

MN8RsHOE00COkRsC#CCDO)0_m
v;
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#ICRF3s	obCMNNO	oNC3D
D;
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0Rv)mR
H#SMoCCOsHRS5
SNSVl$HDR#:R0MsHo=R:RM"N$
";SISSHE80RH:RMo0CC:sR=;Rc
SSSNs88I0H8ERR:HCM0oRCs:(=R;S
SSIDFNs88RH:RMo0CC:sR=;Rj
SSSEEHoNs88RH:RMo0CC:sR=UR(;S
SSL0ND:CRRlsF0DNLCS;
SVS8D:0RRlsFI8Fs
;S2
FSbs50R
SSSq)77RH:RM0R#8F_Do_HOP0COF5sRNs88I0H8ERR-4FR8IFM0R;j2
SSS7amzRF:Rk#0R0D8_FOoH_OPC0RFs58IH0-ERR84RF0IMF2Rj
2SS;S

Ns00H0LkC3R\s	NM\RR:HCM0o;Cs
RRRR0N0skHL0\CR3lsCF_PCMIF_N\sMRH:RMo0CC
s;CRM8CHM00)$Rm
v;
ONsECH0Os0kCCR#D0CO_v)mRRFV)RmvHS#
ObFlFMMC0mR)vN_L#SC
SMoCCOsHRS5
SISSHE80RH:RMo0CC
s;SSSSNs88I0H8ERR:HCM0o;Cs
SSSSIDFNs88RH:RMo0CC
s;SSSSEEHoNs88RH:RMo0CC
s;SSSS0DNLCRR:s0FlNCLD;S
SSVS8D:0RRlsFI8Fs
2SS;S
Sb0FsRS5
SqSS7R7):MRHR8#0_oDFHPO_CFO0sNR58I8sHE80R4-RRI8FMR0Fj
2;SSSS7amzRF:Rk#0R0D8_FOoH_OPC0RFs58IH0-ERR84RF0IMF2Rj
SSS2S;
CRM8ObFlFMMC0
;
SMOF#M0N00RMLRR:HCM0oRCs:4=Rn
;
SMVkOF0HM0R#N)s0FHlpMsCRCs0kMMRH0CCos#RH
PSSNNsHLRDC#CHxRH:RMo0CC
s;SFSOMN#0ML0RD	FO#CHxRH:RMo0CC:sR=0RMLRR*n
c;SoLCHSM
SRHV5IDFNs88R8lFRFLDOH	#xRC2=jRRRC0EMS
SS0sCkRsMDNFI8R8s+DRLF#O	H;xC
CSSD
#CSsSSCs0kM5R5DNFI8R8s+DRLF#O	HRxC-2R4RL/RD	FO#CHx2RR*LODF	x#HCS;
S8CMR;HV
MSC8kRVMHO0F#MR00Ns)pFlH;MC
O
SF0M#NRM0LODF	x#HCRR:HCM0oRCs:n=RcRR*M;0L
FSOMN#0MD0RH8lq8:sRR0HMCsoCRR:=#s0N0l)FpCHM;SR
O#FM00NMR_MLs_FlVOsNRH:RMo0CC:sR=ER5HNoE8R8s-HRDl8q8sRR+4R2/LODF	x#HCS;
O#FM00NMRVDC0F_sls_VN:ORR0HMCsoCRR:=5oEHE8N8sRR-DqHl8R8s+2R4R8lFRFLDOH	#x
C;
$S0b0CRNCLD_k8F0#RHRsNsN5$RMsL_FVl_s+NO4FR8IFM0RRj2FsVRFFlIs
8;
HS#oDMNRk8F0F_slRR:0DNLCF_8k
0;LHCoMS

HLV_Hmo)vH:RVER5HNoE8R8s-FRDI8N8sRR+4RR>LODF	x#HCo2RCsMCN
0CSHS#oDMNRk8F0H_Vs,#0Rz7mak_NGRR:sIFlF;s8
#SSHNoMD7Rq7N)_kRG,q)77_:VRR8#0_oDFHPO_CFO0sNR58I8sHE80R4-RRI8FMR0Fj
2;SoLCH
M
SFSVsH_bbRC:VRFsHMRHR0jRF8RN8HsI8-0E4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#jS;
S0SN0LsHkR0C\N3sMR	\FsVRCAo#RD:RNDLCRRH#4R;
RRRRRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;R
RRRRRRRRRR0RN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
LSSCMoH
SSSs#Coqb:RHLbCkSV
SFSbsl0RN
b5SSSSSRRQ=q>R757)H
2,SSSSRmSRRR=>q)77_HV52S
SS2SS;S

SCSso:#ARbbHCVLk
SSSb0FsRblN5S
SSRSSQ>R=R7q7)5_VH
2,SSSSRmSRRR=>q)77_GNk5
H2SSSSS
2;SMSC8CRoMNCs0VCRFbs_H;bC
S
S) mv4:(RRv)m_#LNCS
SSMoCCOsHRblN5S
SSHSI8R0ES>S=R8IH0
E,SSSSNs88I0H8ESRR=N>R8I8sHE80,SR
SDSSF8IN8RsRR>S=RIDFNs88,S
SSHSEo8EN8RsRR>S=RlDHqs88-
4,SSSS0DNLCRRRSR=>0DNLCS,
S8SSVRD0RSRS=8>RV
D0S2SS
SSSb0FsRblNRR5Rq)77RR=>q)77_RV,
SSSS7SSmRza=8>RF_k0V#Hs0S
SS2SS;
S
SFS8ks0_Fjl52=R<Rk8F0H_VsR#0IMECR75q7N)_k>GR=mRBh1e_ap7_mBtQ_Be a5m)DNFI8,8sR8N8s8IH02E2
SSSSSSSSRRRCCD#RD8V0
;
SFSVsF_DFRb:VRFsHMRHR04RFLRM_lsF_NVsOCRoMNCs0SC
SHS#oDMNRk8F00_#NRoC:FRslsIF8S;
SoLCHSM
SmS)vR 6:mR)vN_L#SC
SCSoMHCsONRlbS5
SISSHE80R=SS>HRI8,0E
SSSS8N8s8IH0RERSR=>Ns88I0H8E
,RSSSSDNFI8R8sR=RS>HRDl8q8sRR+54H-2D*LF#O	H,xC
SSSSoEHE8N8sRRRSR=>DqHl8R8s+*RHLODF	x#HC,-4RS
SSNS0LRDCR=RS>NR0L,DC
SSSSD8V0RRRS>S=RD8V0S
SSS2
SFSbsl0RN5bRR7Rq7=)R>7Rq7V)_,SR
SSSSSz7ma>R=Rk8F00_#N
oCSSSSSS2;
S
SSk8F0F_sl25HRR<=80Fk_N#0oICRERCM57q7)k_NG=R>RhBmea_17m_pt_QBea BmD)5H8lq85s+H2-4*FLDOH	#xRC,Ns88I0H8E
22SSSSSSSSRCRRDR#C80Fk_lsF54H-2S;
S8CMRMoCC0sNCFRVsF_DF
b;SS
SH#V_H:xCRRHV5VDC0F_sls_VN>ORRRj2oCCMsCN0
SSS#MHoN8DRF_k0#o0NCRR:sIFlF;s8
LSSCMoH
SSS) mv6RR:)_mvLCN#
SSSoCCMsRHOl5Nb
SSSS8IH0SERSR=>I0H8ES,
SNSS8I8sHE80R=RS>8RN8HsI8,0ERS
SSFSDI8N8sRRRSR=>DqHl8R8s+LRM_lsF_NVsOD*LF#O	H,xC
SSSSoEHE8N8sRRRSR=>EEHoNs88,SR
S0SSNCLDRSRR=0>RNCLD,S
SSVS8DR0RR=SS>VR8DS0
S
S2SbSSFRs0lRNb5qRR7R7)=q>R7_7)V
,RSSSSSmS7z=aR>FR8k#0_0CNo
SSSS;S2S

SS8SSF_k0s5FlMsL_FVl_s+NO4<2R=FR8ks0_FMl5LF_sls_VN
O2SSSSSSSSSISSERCM57q7)k_NGRR<Bemh_71a_tpmQeB_ mBa)H5Dl8q8sL+M_lsF_NVsOD*LF#O	H,xCR8N8s8IH02E2
SSSSSSSSRRRSRSRRDRC#8CRF_k0#o0NCS;

SSS7amz_GNkRR<=80VDRCIEMqR57_7)NRkG>mRBh1e_ap7_mBtQ_Be a5m)EEHoNs88,8RN8HsI820E2S
SSSSSSDRC#8CRF_k0s5FlMsL_FVl_s+NO4
2;SMSC8CRoMNCs0HCRVH_#x
C;SS
SHMV_#CHx:VRHRC5DVs0_FVl_sRNO=2RjRMoCC0sNCS
SSz7mak_NG=R<RD8V0ERIC5MRq)77_GNkRB>Rm_he1_a7pQmtB _eB)am5oEHE8N8sN,R8I8sHE802S2
SSSSSCSRDR#C80Fk_lsF5_MLs_FlVOsN2S;
S8CMRMoCC0sNCVRH_HM#x
C;
VSSFbs_H:bCRsVFRHHRMRRj0IFRHE80-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#.R;
RRRRRRRRRNRR0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RSSLHCoMS
SSCRsoR#:bCHbL
kVSSSSRsbF0NRlbS5
SRRRSSSSRRRQ=7>Rm_zaN5kGH
2,SRSRRSSSSmRRRR=>7amz5
H2SSSSS2SR;S
SR8CMRMoCC0sNCFRVsH_bb
C;
MSC8CRoMNCs0HCRVH_Lov)m;S

H#V_lDND):mvRRHV5oEHE8N8sRR-DNFI8R8s+RR4<L=RD	FO#CHx2CRoMNCs0SC
So#HMRNDq)77_:VRR8#0_oDFHPO_CFO0sNR58I8sHE80R4-RRI8FMR0Fj
2;SoLCHSM
SsVF_bbHCV:RFHsRRRHMjFR0R8N8s8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;S
SLHCoMS
SSosC#Rq:bCHbL
kVSSSSb0FsRblN5S
SSQSSRR=>q)775,H2
SSSSRSm=q>R7_7)V25H
SSSS
2;SMSC8CRoMNCs0VCRFbs_H;bC
)
Sm6v R):RmLv_N
#CSSSSoCCMsRHOl5Nb
SSSSSSSI0H8ESRS=I>RHE80,R
RSSSSSNSS8I8sHE80R=RR>8RN8HsI8,0ERS
SSSSSSIDFNs88RSRR=D>RF8IN8
s,SSSSSESSHNoE8R8sR=RS>HREo8EN8
s,SSSSS0SSNCLDRSRR=0>RNCLD,S
SSSSSSD8V0RRRS>S=RD8V0S
SSSSSSS2
SbSSFRs0lRNb5qRR7R7)=q>R7_7)V
,RSSSSS7SSmRza=7>Rm
zaSSSSS;S2SS

CRM8oCCMsCN0R_HV#DlNDv)m;C

MN8RsHOE00COkRsC#CCDO)0_m
v;
