@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)am_h ]"ma;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"
RHR`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCR
R`8CMH
V
`8HVCmVReqp_1)1 ah_m
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RbRRsCFbsR0$q 11)ma_h] _mXa_Z;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR55!fkH#MF	MI0M5C_#0CsGb2;22
RRRR8CMbbsFC$s0
`RRCHM8V/R/Rpme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RbbsFC$s0R1q1 _)am_h ]_mauR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
Rf!5HM#k	IMFMC50#C0_G2bs2-R|>fR5FEMCF005C_#0CsGb2
2;RMRC8Fbsb0Cs$R

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)am_h ]_mauR:RR#RN#0CsRFbsb0Cs$qR51)1 ah_m m_]a2_u
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HMFROMH0NMl#RFRsCFDsRCR##0MENRN4R#s#C0RC8L#H0"
2;`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 ah_m m_]aZ_X_Ru:NC##sb0RsCFbsR0$51q1 _)am_h ]_maXuZ_2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRR//m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/eRmpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eqp_1v1z RR:LHCoMRR:F_PDNk##lRC
RRRRRvRR_1q1 _)am_h ]_mauR:RR#RN#CklRFbsb0Cs$qR51)1 ah_m m_]a2_u;`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )_ mh_a]m__XZuN:R#l#kCsRbFsbC05$Rq 11)ma_h] _mXa_Z2_u;R
R`8CMH/VR/eRmpv_QuBpQQXa_BB] iw_mwC
`MV8HRR//m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"R2;RRR
RCRRMN8O#
C
RMRC8MoCC0sNC`

CHM8V/R/Rpme_1q1 _)am
h
`8HVCmVReBp_m)e _
mh
RRRRIRRHRsCr8IH04E-:Rj900C#_bCGsR_4=CR0#C0_GRbs-{R{I0H8E{-44j'L}4},'}L4;R
RRRRRsRCor8IH04E-:Rj9F_MCE#F0_COEO8	C;

RRCRoMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )1QqhamY_hL2RCMoHRF:RPOD_FsPC_M#NH
0$
RRRRORRFsPC_#0C0G_CbOs_EoNMCR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R`55m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRfR!#L0ND0C5C_#0CsGb22R2
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_NOEMRoCOCFPs"C82R;
RRRRCRM8/N/#M$H0RPOFCosNCR

RRRRH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR

RRRRRINDNR$#@b@5F8#CoOCRDR	2LHCoMR
RRRRRRVRHRm5`e)p_ a1 _t1QhRqp!4=R'2LjRoLCHRM
RRRRRRRRRRHV5C50#C0_GRbs^CR0#C0_G2bs=I={HE80{L4'j2}}RoLCHRM
RRRRRRRRRHRRV!R55C50#C0_GRbs={=RI0H8E'{4L}j}2|R|
RRRRRRRRRRRRRRRR5RR00C#_bCGsRR&00C#_bCGs2_4RR!={8IH04E{'}Lj}R22LHCoMR
RRRRRRRRRRRRRF_MCE#F0_COEO8	CRR<=F_MCE#F0_COEO8	CR0|RC_#0CsGb;R
RRRRRRRRRRMRC8R
RRRRRRRRRC
M8RRRRRRRRC
M8RRRRRRRRCCD#RoLCH`M
HCV8VeRmph_QQ)a_ Rt
RRRRRRRRF_MCE#F0_COEO8	CRR<={8IH04E{'}Lj}`;
CHM8VR
RRRRRRMRC8RRRRRRRR
RRRRRRRMRC8/R/RINDN
$#
RRRRORRFsPC_DND_CFM_0EF#E_OCCO	8R:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	RFfs#FC5MEC_F_0#OOEC	RC8={=RI0H8E'{4L}4}2R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"DND_CFM_0EF#E_OCCO	8FROPCCs8;"2
R
RRCRRM/8R/sOFMRCsOCFPsCNo
RRRR8CM
R
RCoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
