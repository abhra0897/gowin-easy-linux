`ifndef ATCMSTMUX100_CONST_VH
`define ATCMSTMUX100_CONST_VH

`define	ATCMSTMUX100_PRODUCT_ID	32'h000c1002

`endif
