-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRR:1RR08NMNRs8ep]7RM1$0#ECHu#RNNO	o
C#-R-RRRRRRRRRR:RRRhR5z)v Q1B_az7_ht1QhR 7b	NONRoC8DCON0sNH2FM
R--RRRRRRRRRRRR:-
-RpRRHNLssR$RRR:Ra#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRRR:R#L$lFODHN$DDRlMNCQ8R 3  
R--RRRRRRRRRRRR:-
-R7RRCDPCFsbC#R:RqCOODsDCN]Re7ap-BN,RMQ8R R  u(4jnFRWsM	HosRtF
kb-R-RRRRRRRRRR:RR
R--RkRus#bFCRRR:aRRERH#b	NONRoC8HCVMRC#MCklsRHO0C$b#MRN8sRNHl0ECO0HRMVkOF0HM-#
-RRRRRRRRRRRRRR:RsVFRCk#R0IHE$R#MC0E#RH#0DFF#e3RNCDk#VRFRb0$CaR17p_zmBtQ_Be a
m)-R-RRRRRRRRRR:RRRsRNCMRH0bCssCC08#RNR#kMHCoM8kRMlsLC#MRHROPC0RFsVlFs3-
-RRRRRRRRRRRRRR:RaRECD0CVl0F#R0LHRRH#0NsC0RC8N0#RElCRFR#0#MHoHOVHNRM0L3H0
R--RRRRRRRRRRRR:aRRERH#b	NONRoCO0FMN#HMRCFPsNDF8RC8N0sHE0lCHFORbNCs0#FsR
FM-R-RRRRRRRRRR:RRRER0CaR17p_zmBtQ_Be aRm)0C$b3ERaCNRbOo	NCDRN#OFRFNM0H
M#-R-RRRRRRRRRR:RRR#RkCDVkRb0$CFROMsPC#MHF#kRVMHO0F,M#RFODO8	RCO0C0MHF
R--RRRRRRRRRRRR:VRRk0MOH#FM,MRN80RFERCskD0HHR0$VOkM0MHF#-3
-RRRRRRRRRRRR
R:-R-RRRRRRRRRR:RRRVRQR$NMRoNskMlC0FR0RVNRk0MOHRFMHN#RRDMkDsRNs,N$RMNRkRDDNNss$-
-RRRRRRRRRRRRRR:RHs#RCs0kMRC85OCGCHb0F,M#RRHVN,M$RCNsR0MFCH8RMP8HHN8kD2D$3-
-
R--RFRh0RCRRRRR:aRRERH#b	NONRoClRN$LlCRFV8HHRC80HFRMkOD8NCR808HHNFMDNR80-N
-RRRRRRRRRRRRRR:RJsCkCHs8$RLRF0FDR#,LRk0Hl0RkR#0HMMRFNRI$ERONCMoRC0E
R--RRRRRRRRRRRR:CRRGs0CMRNDHCM0sOVNCF#RsHR#lNkD0MHFRELCNFPHsVRFRC0E
R--RRRRRRRRRRRR:8RRCs#OHHb0FRM3QH0R#CRbs#lH#DHLCFR0R8N8RlOFl0CM#MRN8s/F
R--RRRRRRRRRRRR:NRR0H0sLCk0#FR0RC0ERObN	CNoRO8CDNNs0MHF#L,RkM0RF00RFERONCMo
R--RRRRRRRRRRRR:FRRsCR8DCC0R$NMRHFsoNHMDHRDMRC#F0VREbCRNNO	o8CRCNODsHN0F
M3-R-RRRRRRRRRR:RRRERaCNRbOo	NCFRL8l$RNL$RCERONCMo8MRFDH$RMORNO8FsNCMOR0IHE-
-RRRRRRRRRRRRRR:R0REC0lCs#VRFRNBDkR#C4FnRVER0H##R08NMN3s8
R--RRRRRRRRRRRR:-
-R---------------------------------------------------------------------
-RCf)PHH#FRM:4j..R-f
-7RfN:0CRj.jUc-j-R4j44(:ng:jRg+jd5jRa,EkRR4jqRbs.Ujj2
Rf---R-----------------------------------------------------------------
--
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;b	NONRoCh zv)_QB1_a7zQh1t7h R
H#RFROMN#0MB0RF)b$H0oEhHF0O:CRR)1aQRht:R=
R"RRB$FbsEHo0jR.jQUR 3  RDqDRosHER0#sCC#s8PC3
";
-RR-8RQ:3RqdR
RVOkM0MHFR""+R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5XvqQvvz5pp' aht]),R'hp t2a]-84RF0IMF2Rj3R
R-)-RCD#k0q:R8R8#0RIFzQh1t7h ROPC0#FsRN0E0NRl$CRLRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8Rdq3)R
RVOkM0MHFR""+5:pRR71a_mzpt_QBea BmR);)RR:1_a7ztpmQRB2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5pp' aht]R-48MFI0jFR2R
R-)-RCD#k01:RHDlHN0sRF3RqdERICRsC)#RHRFNRMLCRH10Raz7_pQmtB _eB)am
R
R-Q-R8q:R3
dpRkRVMHO0F"MR+p"5R1:Raz7_pQmtB);RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea Bm))5'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Rl1HHsDNRR0FqR3dIsECCRRpHN#RRCFMR0LHR1zhQ th7R

RR--QR8:q
36RkRVMHO0F"MR+5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5pp' aht]R-48MFI0jFR2R3
RR--)kC#DR0:q#88RRNMzQh1t7h ROPC0,FsRRp,IEH0RMNRFMM-C0oNHRPCQ hat, )R
)3
-RR-8RQ:3RqnR
RVOkM0MHFR""+RR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea Bm))5'hp t-a]4FR8IFM0R3j2
-RR-CR)#0kD:8Rq8N#RRMMF-oMCNP0HChRQa  t)p,R,HRI0NERMhRz1hQt P7RCFO0s),R3R

R=--=========================================================================
==
-RR-8RQ:3RqgR
RVOkM0MHFR""-R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7vQqXv5zvp 'ph]ta,'R)pt ha-]24FR8IFM0R3j2
-RR-CR)#0kD:kR1LN0sOR0#0RIFzQh1t7h ROPC0#FsRN0E0NRl$CRLRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8Rgq3)R
RVOkM0MHFR""-5:pRR71a_mzpt_QBea BmR);)RR:1_a7ztpmQRB2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5pp' aht]R-48MFI0jFR2R
R-)-RCD#k01:RHDlHN0sRF3RqgERICRsC)#RHRFNRMLCRHz0Rht1Qh
 7
-RR-8RQ:3RqgRp
RMVkOF0HM-R""R5p:aR17p_zmBtQ;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQeB_ mBa)'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1HHlDRNs0qFR3IgRECCsRHpR#RRNFRMCLRH0zQh1t7h 
R
R-Q-R8q:R3
44RkRVMHO0F"MR-5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5pp' aht]R-48MFI0jFR2R3
RR--)kC#DR0:10kLs0NO#RRNM-FMMNCo0CHPRaQh )t ,,R)RFVslMRNR1zhQ th7CRPOs0F,3Rp
R
R-Q-R8q:R3
4.RkRVMHO0F"MR-5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5p)' aht]R-48MFI0jFR2R3
RR--)kC#DR0:10kLs0NO#MRNR1zhQ th7CRPOs0F,,R)RFVslRRNM-FMMNCo0CHPRaQh )t ,3Rp
R
R-=-==========================================================================
=
R-R-R:Q8R4q36R
RVOkM0MHFR""*R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5'5ppt ha)]+'hp t-a]482RF0IMF2Rj3R
R-)-RCD#k0u:RCFsVsRl#0RECl0kDHHbDOHN0FFMRbNCs0MHFRRFM0RIFzQh1t7h ROPC0#Fs
-RR-RRRRRRRRER0Nl0RNb$RFH##LRD$LFCRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8q:R3
4(RkRVMHO0F"MR*5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5'5ppt hap]+'hp t-a]482RF0IMF2Rj3R
R-)-RCD#k0v:RkHD0bCDH#MRNR1zhQ th7CRPOs0F,,RpR0IHERRNM-FMMNCo0CHP
-RR-RRRRRRRRhRQa  t)),R3RR)HO#RFCMPs80CRR0FNzMRht1QhR 7P0COFFsRVR
R-R-RRRRRR1RRQRZ p 'ph]taRVLCFRsCl0kDHHbDOHN0F
M3
-RR-8RQ:3Rq4RU
RMVkOF0HM*R""pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)5p)' aht]'+)pt ha4]-2FR8IFM0R3j2
-RR-CR)#0kD:kRvDb0HD#HCRRNMzQh1t7h ROPC0,FsRR),IEH0RMNRFMM-C0oNH
PCR-R-RRRRRRRRRaQh )t ,3RpRHpR#FROMsPC0RC80NFRMhRz1hQt P7RCFO0sVRF
-RR-RRRRRRRRQR1Z) R'hp tRa]LFCVslCRkHD0bODHNF0HM
3
R-R-============================================================================
-RR-R
R-h-Rm:a RRQV#FCOMN8RslokCRM0Hx#RCRsFVRFs"R/"FsbCNs0F,RRN#CCPs$H0RPDCCRD
RR--RRRRRVRFR) )mH)R##RH#8kC3R

RR--QR8:q43.
VRRk0MOHRFM"R/"5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#MRNR1zhQ th7CRPOs0F,,RpRRL$N0MFERCszQh1t7h ROPC0,FsR
)3
-RR-8RQ:3Rq.Rd
RMVkOF0HM/R""pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#MRNR1zhQ th7CRPOs0F,,RpRRL$NFRMMC-MoHN0PQCRhta  R),)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:qc3.
VRRk0MOHRFM"R/"5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQeB_ mBa)'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#NFRMMC-MoHN0PQCRhta  R),pL,R$MRNR1zhQ th7CRPOs0F,3R)
-RR-RRRRRRRRVRQR_hmmAw_Q5a1p>2RRp)' aht]s,RCD#k0#RHRk0sM0ONC08RF'R)pt ha
]3
-RR-============================================================================R
R-R-
RR--h ma:VRQRO#CFRM8Nksol0CMRRH#xFCsRsVFRC"slF"RbNCs0,FsR#NRCsPCHR0$DCCPDR
R-R-RRRRRRRFV m)))#RHR#H#k3C8
R
R-Q-R8q:R3
.(RkRVMHO0F"MRs"ClR,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5p)' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#Fs3R

RR--QR8:qg3.
VRRk0MOHRFM"lsC"pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpCRsl"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRM)8RRRH#NR
R-R-RRRRRRMRRFMM-C0oNHRPCQ hat3 )
-RR-RRRRRRRRVRQR_hmmAw_Q5a1)>2RRpp' aht]s,RCD#k0#RHRk0sM0ONC08RF'Rppt ha
]3
-RR-8RQ:3RqdRj
RMVkOF0HMsR"CRl"5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQeB_ mBa)'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRH)R#MRNR1zhQ th7CRPOs0FR8NMRHpR#
RNR-R-RRRRRRRRRMMF-oMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0F) 'ph]ta3R

R=--=========================================================================
==R-R-
-RR-mRhaR :Q#VRCMOF8sRNoCklMH0R#CRxsVFRF"sRl"F8RCFbsFN0sN,RRP#CC0sH$CRDP
CDR-R-RRRRRFRRV)R )Rm)HH#R#C#k8
3
R-R-R:Q8Rdq3dR
RVOkM0MHFRF"l85"Rp),RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea Bm))5'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"R8lFRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0s
#3
-RR-8RQ:3RqdR6
RMVkOF0HMlR"FR8"5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsM1_a7ztpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQeB_ mBa)'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"plRF8)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NMRR)
RR--RRRRRRRRHN#RRMMF-oMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:qn3d
VRRk0MOHRFM"8lF"pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpFRl8"R)RCIEs)CRRRH#NzMRht1QhR 7P0COFNsRMp8R
-RR-RRRRRRRR#RHRMNRFMM-C0oNHRPCQ hat3 )
-RR-RRRRRRRRVRQR_hmmAw_Q5a1p>2RRp)' aht]s,RCD#k0#RHRk0sM0ONC08RF'R)pt ha
]3
-RR-============================================================================R
R-Q-R8q:R3
dgRkRVMHO0FVMRH_M8D0CVl0F#R)5qtRR:1_a7ztpmQeB_ mBa)Y;RR1:Raz7_pQmtBs2RCs0kMhRQa  t)R;
RR--)kC#D#0Rk$L0bRC:Q hat
 )R-R-R#)Ck:D0RMwH80#REDCRClV0FR#0FkOOsMsCOFCRVER0CNRPDRkCFYVRRRHMq3)t
-RR-RRRRRRRRCR)0Mks#ER0CMRH8RCGF0VREFCROsOksOCMCVRHRRH0C#GH0R#,F-sR40RFEICsH3#C
R
R-Q-R8q:R3
c4RkRVMHO0FVMRH_M8sEHo0#lF0qR5):tRR71a_mzpt_QBea BmR);YRR:1_a7ztpmQRB2skC0sQMRhta  
);R-R-R#)CkRD0#0kL$:bCRaQh )t 
-RR-CR)#0kD:HRwMR8#0RECD0CVl0F#ROFOkCssMROCF0VREPCRNCDkRRFVYMRHRtq)3R
R-R-RRRRRR)RRCs0kM0#REHCRMG8CRRFV0RECFkOOsMsCOHCRV0RHRHCG#,0#RRFs-F4R0sECICH#3R

R=--=========================================================================
==R-R-RlBFbHNs#RFMmsbCNs0F#R
R-=-==========================================================================
=
R-R-R:Q8R4B3
VRRk0MOHRFM"R>"5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3Rd
RMVkOF0HM>R""pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCp#RHRMNRFMM-C0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:B
36RkRVMHO0F"MR>5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMF-oMCNP0HChRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3R(
RMVkOF0HM<R""pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RgB3
VRRk0MOHRFM"R<"5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB4R4
RMVkOF0HM<R""pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNM-FMMNCo0CHPRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RB4Rd
RMVkOF0HM<R"=5"Rp),RR1:Raz7_pQmtB _eB)am2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
46RkRVMHO0F"MR<R="5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NFRMMC-MoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
4(RkRVMHO0F"MR<R="5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R4B3gR
RVOkM0MHFR=">"pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB.R4
RMVkOF0HM>R"=5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB.Rd
RMVkOF0HM>R"=5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMC-MoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:B63.
VRRk0MOHRFM"R="5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
.(RkRVMHO0F"MR=5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRHpR#RRNM-FMMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8R.B3gR
RVOkM0MHFR""=RR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8RdB34R
RVOkM0MHFR="/"pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBdRd
RMVkOF0HM/R"=5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBdR6
RMVkOF0HM/R"=5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMC-MoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:B(3d
VRRk0MOHRFMvQQhvRzv5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a
m)R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsF0VRIzFRht1QhR 7P0COFRs#00ENR$lNR
LCR-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RdB3gR
RVOkM0MHFRhvQQvvzRR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea BmR)
RR--)kC#DR0:)kC0sRM#0RECD#C#CFsRVRRNMMFMC0oNHRPCQ hat, )RRp,N
M8R-R-RRRRRRRRRRNMzQh1t7h ROPC0,FsR
)3
-RR-8RQ:3RBcR4
RMVkOF0HMQRvhzQvvpR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a
m)R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRMhRz1hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRRMMFMNCo0CHPRaQh )t ,3R)
R
R-=-==========================================================================
=
R-R-R:Q8RcB3dR
RVOkM0MHFRXvqQvvzR,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am
-RR-CR)#0kD:CR)0Mks#ER0CsRoCCN0sVRFRF0IR1zhQ th7CRPOs0F#ER0Nl0RNL$RCR
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
c6RkRVMHO0FvMRqvXQz5vRpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am
-RR-CR)#0kD:CR)0Mks#ER0CsRoCCN0sVRFRMNRFCMMoHN0PQCRhta  R),pN,RMR8
RR--RRRRRRRRNzMRht1QhR 7P0COFRs,)
3
R-R-R:Q8RcB3(R
RVOkM0MHFRXvqQvvzRR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea BmR)
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsFNVRMhRz1hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRRMMFMNCo0CHPRaQh )t ,3R)
R
R-=-==========================================================================R=
RR--QR8:Bg3c
VRRk0MOHRFM""?>R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB6R4
RMVkOF0HM?R">5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB6Rd
RMVkOF0HM?R">5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:B636
VRRk0MOHRFM""?<R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB6R(
RMVkOF0HM?R"<5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB6Rg
RMVkOF0HM?R"<5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:B43n
VRRk0MOHRFM"=?<"pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bd3n
VRRk0MOHRFM"=?<"pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBnR6
RMVkOF0HM?R"<R="5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RBnR(
RMVkOF0HM?R">R="5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBnRg
RMVkOF0HM?R">R="5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:B43(
VRRk0MOHRFM"=?>"pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:Bd3(
VRRk0MOHRFM""?=R,5pR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB(R6
RMVkOF0HM?R"=5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB(R(
RMVkOF0HM?R"=5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-============================================================================R

RR--QR8:Bg3(
VRRk0MOHRFM"=?/"pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B43U
VRRk0MOHRFM"=?/"pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBURd
RMVkOF0HM?R"/R="5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

R=--=========================================================================
==R-R-RH1EVN0RM)8RF00NCkRwMHO0F
M#R-R-============================================================================
R
R-Q-R81:R3R4
RMVkOF0HM]R1Q_wapa wR)5qtRR:1_a7ztpmQeB_ mBa)B;RmazhRh:Rq)azq
p2RRRRskC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRN#VEH0C-DVF0RMMRNR1zhQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0R''j3R
R-R-RRRRRRaRREBCRmazhRVDC0#lF0DRCCMlC0N#RsDCRF3#0
R
R-Q-R81:R3R.
RMVkOF0HM]R1Q_wa)]QtaqR5):tRR71a_mzpt_QBea BmR);BhmzaRR:hzqa)2qp
RRRR0sCkRsM1_a7ztpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRN#VEH0H-soRE0FNMRMhRz1hQt P7RCFO0smRBzRha0CHl#R3
RR--RRRRRRRRaRECPNNO0RC8bHF#0MHF#sRNCHRVD8DCR0IHEjR''R3
RR--RRRRRRRRaRECBhmzaHRsolE0FR#0ClDCC#M0RCNsR#DF0R3
R=--=========================================================================
==
-RR-8RQ:3R16R
RVOkM0MHFRa)mq_a pa wR)5qtRR:1_a7ztpmQeB_ mBa)B;RmazhRh:Rq)azq
p2RRRRskC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRNsNF00DC-CRV0FNVRMhRz1hQt P7RCFO0smRBzRha0CHl#
3
R-R-R:Q8Rn13
VRRk0MOHRFM)qmaa) _Qat]R)5qtRR:1_a7ztpmQeB_ mBa)B;RmazhRh:Rq)azq
p2RRRRskC0s1MRaz7_pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB _eB)am5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRNsNF00sC-H0oERRFVNzMRht1QhR 7P0COFBsRmazhRl0HC
#3
R
R-=-==========================================================================
=
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413(#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14R(
RMVkOF0HM#R"DRN"5tq)R1:Raz7_pQmtB _eB)am;mRBzRha:hRQa  t)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]Qa _pwqa5)Rt,Bhmza
2
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413g#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14Rg
RMVkOF0HM#R"sRN"5tq)R1:Raz7_pQmtB _eB)am;mRBzRha:hRQa  t)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be a5m)q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]QaQ_)t5]aq,)tRzBmh
a2
R
R-=-==========================================================================R=
RR--R R)1 QZRMwkOF0HMR#
R=--=========================================================================
==
-RR-8RQ:3R).R
RVOkM0MHFR1) QRZ 5tq)R1:Raz7_pQmtB _eB)am; RhWQ_1Z: RRahqzp)q2R
RRCRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea Bmh)5 1W_Q-Z 4FR8IFM0R
j2R-R-R#)Ck:D0R#)CH#xCRC0ER1zhQ th7CRPOs0FRtq)RR0F0REC#ObCHCVH8HR#x
C3R-R-RRRRRRRRRRaFONsC0NCRRsDNoRCsP0COFRs,0RECMRCIrVDC0#lF0L9RHb0RF0#HH#FM
-RR-RRRRRRRRsRNCHRVD8DCR0IHEjR''W3RERCM0MskOHN0MRo,0RECD0CVl0F#R0LH#R
R-R-RRRRRRNRRs8CRsbFbC
83
VRRk0MOHRFM)Q 1Z5 Rq,)tRZ1Q  _)1RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be a;m)
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ_Be aRm)5Z1Q  _)1C'DMEo0-84RF0IMF2Rj
R
R-=-==========================================================================R=
RR--BPFMCHs#FwMRk0MOH#FM
-RR-============================================================================R

RR--QR8:7
34RkRVMHO0FaMRmh_Qa  t)qR5):tRR71a_mzpt_QBea BmR)2skC0shMRq)azq
p;R-R-R#)CkRD0#0kL$:bCRahqzp)q3NReDRkCOMNMFL0RCCRMoHN0P#CRHCMORsbNN0lCCHsR#MRN
-RR-RRRRRRRRRRRRhRz1hQt P7RCFO0sR3
RR--)kC#DR0:BPFMC#s0RC0ER1zhQ th7CRPOs0FRR0FNQMRhta  
)3
-RR-8RQ:3R7dR
RVOkM0MHFR_aF1p08FOoHe0COF5sRq,)tRZ1Q RR:hzqa)2qpR0sCkRsM1_a7pQmtB _eB)am;R
R-)-RCD#k0kR#Lb0$C1:Rap7_mBtQ_Be a5m)1 QZ-84RF0IMF2Rj
-RR-CR)#0kD:FRBMsPC0N#RRMMF-oMCNP0HChRQa  t)FR0RRNMzQh1t7h ROPC0RFsIEH0
-RR-RRRRRRRRER0CbR#CVOHHRC81 QZ3R

RMVkOF0HMFRa_810pHFoOOeC0RFs5tq)Rh:Rq)azqRp;1 QZ_1) R1:Raz7_pQmtB _eB)am2R
RRCRs0MksR71a_tpmQeB_ mBa)R;
RR--)kC#D#0Rk$L0bRC:1_a7pQmtB _eB)am5Z1Q  _)1C'DMEo0-84RF0IMF2Rj
R
RNNDH#FRa_810_opFHeO_CFO0s#RH
RRRR_aF1p08FOoHe0COFhsrq)azqRp,hzqa)RqpskC0s1MRap7_mBtQ_Be a9m);R
RNNDH#FRa_e1pR
H#RRRRa1F_0F8poeHOCFO0sqrhaqz)ph,Rq)azqspRCs0kMaR17m_pt_QBea Bm;)9
NRRD#HNR_aF1_08pHFoOC_eOs0FR
H#RRRRa1F_0F8poeHOCFO0sqrhaqz)p1,Raz7_pQmtB _eB)amR0sCkRsM1_a7pQmtB _eB)am9R;
RHNDNa#RFp_1e#RH
RRRR_aF1p08FOoHe0COFhsrq)azqRp,1_a7ztpmQeB_ mBa)CRs0MksR71a_tpmQeB_ mBa)
9;
-RR-8RQ:3R76R
RVOkM0MHFR_aF1z08pHFoOOeC0RFs5tq),QR1Z: RRahqzp)q2CRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_mzpt_QBea Bm1)5Q-Z 4FR8IFM0R
j2R-R-R#)Ck:D0RMBFP0Cs#RRNM-FMMNCo0CHPRaQh )t RR0FNzMRht1QhR 7P0COFIsRH
0ER-R-RRRRRRRRRC0ERC#bOHHVC18RQ3Z 
R
RVOkM0MHFR_aF1z08pHFoOOeC0RFs5tq)Rh:Rq)azqRp;1 QZ_1) R1:Raz7_pQmtB _eB)am2R
RRCRs0MksR71a_mzpt_QBea Bm
);R-R-R#)CkRD0#0kL$:bCR71a_tpmQeB_ mBa)Q51Z) _ D1'C0MoER-48MFI0jFR2R

RHNDNa#RF0_18p_zFOoH_OeC0RFsHR#
RaRRF0_18FzpoeHOCFO0sqrhaqz)ph,Rq)azqspRCs0kMaR17p_zmBtQ_Be a9m);R
RNNDH#FRa_p1ze#RH
RRRR_aF1z08pHFoOOeC0rFshzqa),qpRahqzp)qR0sCkRsM1_a7ztpmQeB_ mBa)
9;RDRNHRN#a1F_0z8_pHFoOC_eOs0FR
H#RRRRa1F_0p8zFOoHe0COFhsrq)azqRp,1_a7ztpmQeB_ mBa)CRs0MksR71a_mzpt_QBea Bm;)9
NRRD#HNR_aF1ezpR
H#RRRRa1F_0p8zFOoHe0COFhsrq)azqRp,1_a7ztpmQeB_ mBa)CRs0MksR71a_mzpt_QBea Bm;)9
M
C8NRbOo	NCzRhvQ )Ba_17h_z1hQt 
7;
LDHs$NsRCHCCk;
#HCRC3CCMCkls_HO#308N;DD
N
bOo	NCFRL8h$Rz)v Q1B_az7_ht1QhR 7H
#
R-R-R:Q8Rdq3
VRRk0MOHRFM"R+"5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)51zhQ th725pRz+Rht1Qh5 7);22
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3
d)RkRVMHO0F"MR+p"5R1:Raz7_pQmtB _eB)am;RR):aR17p_zmBtQ2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RzQh1t7h 5Rp2+2R);R
RCRM8VOkM0MHFR""+;R

RR--QR8:qp3d
VRRk0MOHRFM"5+"pRR:1_a7ztpmQRB;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)5+pRR1zhQ th725)2R;
R8CMRMVkOF0HM+R""
;
R-R-R:Q8R6q3
VRRk0MOHRFM"R+"5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)zR5ht1Qh5 7p+2RR;)2
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3Rn
RMVkOF0HM+R""pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)5+pRR1zhQ th725)2R;
R8CMRMVkOF0HM+R""
;
R-R-============================================================================
R
R-Q-R8q:R3Rg
RMVkOF0HM-R""pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)zR5ht1Qh5 7p-2RR1zhQ th725)2R;
R8CMRMVkOF0HM-R""
;
R-R-R:Q8Rgq3)R
RVOkM0MHFR""-5:pRR71a_mzpt_QBea BmR);)RR:1_a7ztpmQRB2skC0s1MRaz7_pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s1MRaz7_pQmtB _eB)amRh5z1hQt p752RR-)
2;RMRC8kRVMHO0F"MR-
";
-RR-8RQ:3RqgRp
RMVkOF0HM-R""R5p:aR17p_zmBtQ;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)pR5Rz-Rht1Qh5 7);22
CRRMV8Rk0MOHRFM";-"
R
R-Q-R8q:R3
44RkRVMHO0F"MR-5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0s1MRaz7_pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s1MRaz7_pQmtB _eB)amRh5z1hQt p752RR-)
2;RMRC8kRVMHO0F"MR-
";
-RR-8RQ:3Rq4R.
RMVkOF0HM-R""pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)5-pRR1zhQ th725)2R;
R8CMRMVkOF0HM-R""
;
R-R-============================================================================
R
R-Q-R8q:R3
46RkRVMHO0F"MR*5"Rp),RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RzQh1t7h 5Rp2*hRz1hQt )752
2;RMRC8kRVMHO0F"MR*
";
-RR-8RQ:3Rq4R(
RMVkOF0HM*R""pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)51zhQ th725pR)*R2R;
R8CMRMVkOF0HM*R""
;
R-R-R:Q8R4q3UR
RVOkM0MHFR""*RR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RpRR*zQh1t7h 52)2;R
RCRM8VOkM0MHFR""*;R

R=--=========================================================================
==
-RR-8RQ:3Rq.R4
RMVkOF0HM/R""pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)zR5ht1Qh5 7p/2RR1zhQ th725)2R;
R8CMRMVkOF0HM/R""
;
R-R-R:Q8R.q3dR
RVOkM0MHFR""/RR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RzQh1t7h 5Rp2/2R);R
RCRM8VOkM0MHFR""/;R

RR--QR8:qc3.
VRRk0MOHRFM"R/"5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)pR5Rz/Rht1Qh5 7);22
CRRMV8Rk0MOHRFM";/"
R
R-=-==========================================================================
=
R-R-R:Q8R.q3(R
RVOkM0MHFRC"sl5"Rp),RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RzQh1t7h 5Rp2sRClzQh1t7h 52)2;R
RCRM8VOkM0MHFRC"sl
";
-RR-8RQ:3Rq.Rg
RMVkOF0HMsR"CRl"5:pRR71a_mzpt_QBea BmR);)RR:hzqa)2qpR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)zR5ht1Qh5 7ps2RC)lR2R;
R8CMRMVkOF0HMsR"C;l"
R
R-Q-R8q:R3
djRkRVMHO0F"MRs"ClRR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RpCRslhRz1hQt )752
2;RMRC8kRVMHO0F"MRs"Cl;R

R=--=========================================================================
==
-RR-8RQ:3RqdRd
RMVkOF0HMlR"FR8"5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)51zhQ th725pR8lFR1zhQ th725)2R;
R8CMRMVkOF0HMlR"F;8"
R
R-Q-R8q:R3
d6RkRVMHO0F"MRl"F8RR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RzQh1t7h 5Rp2lRF8)
2;RMRC8kRVMHO0F"MRl"F8;R

RR--QR8:qn3d
VRRk0MOHRFM"8lF"pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)5lpRFz8Rht1Qh5 7);22
CRRMV8Rk0MOHRFM"8lF"
;
R-R-============================================================================
-RR-8RQ:3RqdRg
RMVkOF0HMHRVMD8_ClV0FR#05tq):aR17p_zmBtQ_Be a;m)RRY:1_a7ztpmQRB2skC0sQMRhta  H)R#R
RLHCoMR
RRCRs0MksRMVH8C_DVF0l#z05ht1Qh5 7q2)t,2RY;R
RCRM8VOkM0MHFRMVH8C_DVF0l#
0;
-RR-8RQ:3RqcR4
RMVkOF0HMHRVMs8_H0oEl0F#R)5qt1:Raz7_pQmtB _eB)am;:RYR71a_mzpt2QBR0sCkRsMQ hatR )HR#
RoLCHRM
RsRRCs0kMHRVMs8_H0oEl0F#51zhQ th7)5qtR2,Y
2;RMRC8kRVMHO0FVMRH_M8sEHo0#lF0
;
R-R-============================================================================
R
R-Q-R8B:R3R4
RMVkOF0HM>R""pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752RR>zQh1t7h 5;)2
CRRMV8Rk0MOHRFM";>"
R
R-Q-R8B:R3Rd
RMVkOF0HM>R""pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMpRR>zQh1t7h 5;)2
CRRMV8Rk0MOHRFM";>"
R
R-Q-R8B:R3R6
RMVkOF0HM>R""pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2>;R)
CRRMV8Rk0MOHRFM";>"
R
R-=-==========================================================================
=
R-R-R:Q8R(B3
VRRk0MOHRFM"R<"5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2<hRz1hQt )752R;
R8CMRMVkOF0HM<R""
;
R-R-R:Q8RgB3
VRRk0MOHRFM"R<"5:pRRahqzp)q;RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMRRp<hRz1hQt )752R;
R8CMRMVkOF0HM<R""
;
R-R-R:Q8R4B34R
RVOkM0MHFR""<RR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p<2RR
);RMRC8kRVMHO0F"MR<
";
-RR-============================================================================R

RR--QR8:Bd34
VRRk0MOHRFM""<=R,5pR:)RR71a_mzpt_QBea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR<=zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""<=;R

RR--QR8:B634
VRRk0MOHRFM""<=RR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0spMRRR<=zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""<=;R

RR--QR8:B(34
VRRk0MOHRFM""<=RR5p:aR17p_zmBtQ_Be a;m)R:)RRahqzp)q2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p<2R=;R)
CRRMV8Rk0MOHRFM""<=;R

R=--=========================================================================
==
-RR-8RQ:3RB4Rg
RMVkOF0HM>R"=5"Rp),RR1:Raz7_pQmtB _eB)am2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p>2R=hRz1hQt )752R;
R8CMRMVkOF0HM>R"=
";
-RR-8RQ:3RB.R4
RMVkOF0HM>R"=5"RpRR:hzqa);qpR:)RR71a_mzpt_QBea BmR)2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR>pR=hRz1hQt )752R;
R8CMRMVkOF0HM>R"=
";
-RR-8RQ:3RB.Rd
RMVkOF0HM>R"=5"RpRR:1_a7ztpmQeB_ mBa));RRh:Rq)azqRp2skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR>=)R;
R8CMRMVkOF0HM>R"=
";
-RR-============================================================================R

RR--QR8:B63.
VRRk0MOHRFM"R="5Rp,)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2=hRz1hQt )752R;
R8CMRMVkOF0HM=R""
;
R-R-R:Q8R.B3(R
RVOkM0MHFR""=RR5p:qRhaqz)p);RR1:Raz7_pQmtB _eB)am2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0spMRRz=Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR=
";
-RR-8RQ:3RB.Rg
RMVkOF0HM=R""pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2=;R)
CRRMV8Rk0MOHRFM";="
R
R-=-==========================================================================
=
R-R-R:Q8RdB34R
RVOkM0MHFR="/"pR5,RR):aR17p_zmBtQ_Be a2m)R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752=R/R1zhQ th725);R
RCRM8VOkM0MHFR="/"
;
R-R-R:Q8RdB3dR
RVOkM0MHFR="/"pR5Rh:Rq)azqRp;)RR:1_a7ztpmQeB_ mBa)s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMp=R/R1zhQ th725);R
RCRM8VOkM0MHFR="/"
;
R-R-R:Q8RdB36R
RVOkM0MHFR="/"pR5R1:Raz7_pQmtB _eB)am;RR):qRhaqz)ps2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2/)=R;R
RCRM8VOkM0MHFR="/"
;
R-R-============================================================================
R
R-Q-R8B:R3
d(RkRVMHO0FvMRQvhQz5vRp),R:aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)vR5QvhQzzv5ht1Qh5 7pR2,zQh1t7h 52)22R;
R8CMRMVkOF0HMQRvhzQvv
;
R-R-R:Q8RdB3gR
RVOkM0MHFRhvQQvvzR:5pRahqzp)q;:R)R71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s1MRaz7_pQmtB _eB)amRQ5vhzQvv,5pR1zhQ th725)2
2;RMRC8kRVMHO0FvMRQvhQz
v;
-RR-8RQ:3RBcR4
RMVkOF0HMQRvhzQvvpR5:aR17p_zmBtQ_Be a;m)RR):hzqa)2qpR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)vR5QvhQzzv5ht1Qh5 7pR2,);22
CRRMV8Rk0MOHRFMvQQhv;zv
R
R-=-==========================================================================R=
RR--QR8:Bd3c
VRRk0MOHRFMvQqXvRzv5Rp,)1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RvQqXv5zvzQh1t7h 5,p2R1zhQ th725)2
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcR6
RMVkOF0HMqRvXzQvvpR5:qRhaqz)p);R:aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)vR5qvXQzpv5,hRz1hQt )752;22
CRRMV8Rk0MOHRFMvQqXv;zv
R
R-Q-R8B:R3
c(RkRVMHO0FvMRqvXQz5vRp1:Raz7_pQmtB _eB)am;:R)Rahqzp)q2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)RvQqXv5zvzQh1t7h 5,p2R2)2;R
RCRM8VOkM0MHFRXvqQvvz;R

R=--=========================================================================
==
-RR-8RQ:3RBcRg
RMVkOF0HM?R">5"Rp),R:aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?>zQh1t7h 5;)2
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:B436
VRRk0MOHRFM""?>R:5pRahqzp)q;:R)R71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp>R?R1zhQ th725);R
RCRM8VOkM0MHFR>"?"
;
R-R-R:Q8R6B3dR
RVOkM0MHFR>"?"pR5:aR17p_zmBtQ_Be a;m)RR):hzqa)2qpR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR1zhQ th725pRR?>)R;
R8CMRMVkOF0HM?R">
";
-RR-============================================================================R

RR--QR8:B636
VRRk0MOHRFM""?<R,5pRR):1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R<hRz1hQt )752R;
R8CMRMVkOF0HM?R"<
";
-RR-8RQ:3RB6R(
RMVkOF0HM?R"<5"Rph:Rq)azqRp;)1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMRRp?z<Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
6gRkRVMHO0F"MR?R<"5Rp:1_a7ztpmQeB_ mBa));R:qRhaqz)ps2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R<;R)
CRRMV8Rk0MOHRFM""?<;R

R=--=========================================================================
==
-RR-8RQ:3RBnR4
RMVkOF0HM?R"<R="5Rp,)1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752<R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
ndRkRVMHO0F"MR?"<=R:5pRahqzp)q;:R)R71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp<R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
n6RkRVMHO0F"MR?"<=R:5pR71a_mzpt_QBea BmR);)h:Rq)azqRp2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2?R<=)R;
R8CMRMVkOF0HM?R"<;="
R
R-=-==========================================================================
=
R-R-R:Q8RnB3(R
RVOkM0MHFR>"?=5"Rp),R:aR17p_zmBtQ_Be a2m)R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR1zhQ th725pR=?>R1zhQ th725);R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RBnRg
RMVkOF0HM?R">R="5Rp:hzqa);qpRR):1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0spMRR=?>R1zhQ th725);R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RB(R4
RMVkOF0HM?R">R="5Rp:1_a7ztpmQeB_ mBa));R:qRhaqz)ps2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R>)=R;R
RCRM8VOkM0MHFR>"?=
";
-RR-============================================================================R

RR--QR8:Bd3(
VRRk0MOHRFM""?=R,5pRR):1_a7ztpmQeB_ mBa)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R=hRz1hQt )752R;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(R6
RMVkOF0HM?R"=5"Rph:Rq)azqRp;)1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMRRp?z=Rht1Qh5 7)
2;RMRC8kRVMHO0F"MR?;="
R
R-Q-R8B:R3
((RkRVMHO0F"MR?R="5Rp:1_a7ztpmQeB_ mBa));R:qRhaqz)ps2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0szMRht1Qh5 7p?2R=;R)
CRRMV8Rk0MOHRFM""?=;R

R=--=========================================================================
==
-RR-8RQ:3RB(Rg
RMVkOF0HM?R"/R="5Rp,)1:Raz7_pQmtB _eB)am2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMhRz1hQt p752/R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"/;="
R
R-Q-R8B:R3
U4RkRVMHO0F"MR?"/=R:5pRahqzp)q;:R)R71a_mzpt_QBea BmR)2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp/R?=hRz1hQt )752R;
R8CMRMVkOF0HM?R"/;="
R
R-Q-R8B:R3
UdRkRVMHO0F"MR?"/=R:5pR71a_mzpt_QBea BmR);)h:Rq)azqRp2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h 5Rp2?R/=)R;
R8CMRMVkOF0HM?R"/;="
R
R-=-==========================================================================
=
R-R-R:Q8R413
VRRk0MOHRFM1w]Qa _pw5aRqR)t:aR17p_zmBtQ_Be a;m)RzBmh:aRRahqzp)q2R
RRCRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR8#0_oDFHPO_CFO0s1R5]aQw_wp aM5k#MHoCq85),t2RzBmh2a2;R
RCRM8VOkM0MHFRQ1]wpa_ ;wa
R
R-Q-R81:R3R.
RMVkOF0HM]R1Q_wa)]QtaqR5):tRR71a_mzpt_QBea BmR);BhmzaRR:hzqa)2qp
RRRR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM#_08DHFoOC_POs0FR]51Q_wa)]QtaM5k#MHoCq85),t2RzBmh2a2;R
RCRM8VOkM0MHFRQ1]w)a_Qat];R

R=--=========================================================================
==
-RR-8RQ:3R16R
RVOkM0MHFRa)mq_a pa wR)5qtRR:1_a7ztpmQeB_ mBa)B;RmazhRh:Rq)azq
p2RRRRskC0s1MRaz7_pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s#MR0D8_FOoH_OPC0RFs5a)mq_a pa w5#kMHCoM8)5qtR2,Bhmza;22
CRRMV8Rk0MOHRFM)qmaap _ ;wa
R
R-Q-R81:R3Rn
RMVkOF0HMmR)a qa_t)Q]5aRqR)t:aR17p_zmBtQ_Be a;m)RzBmh:aRRahqzp)q2R
RRCRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR8#0_oDFHPO_CFO0s)R5maaq Q_)t5]akHM#o8MC5tq)2B,Rmazh2
2;RMRC8kRVMHO0F)MRmaaq Q_)t;]a
R
R-=-==========================================================================
=
R-R-R:Q8R413(R
RVOkM0MHFRD"#N5"Rq:)tR71a_mzpt_QBea BmR);BhmzaQ:Rhta  
)2RRRRskC0s1MRaz7_pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s1MRaz7_pQmtB _eB)amRh5z1hQt q75)Rt2#RDNBhmza
2;RMRC8kRVMHO0F"MR#"DN;R

RR--QR8:1g34
VRRk0MOHRFM"N#s"qR5)Rt:1_a7ztpmQeB_ mBa)B;Rmazh:hRQa  t)R2
RsRRCs0kMaR17p_zmBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be aRm)51zhQ th7)5qt#2RsBNRmazh2R;
R8CMRMVkOF0HM#R"s;N"
R
R-=-==========================================================================
=
R-R-R:Q8R.)3
VRRk0MOHRFM)Q 1Z5 RqR)t:aR17p_zmBtQ_Be a;m)RWh _Z1Q RR:hzqa)2qp
RRRR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)
R5RRRRR R)1 QZR)5qtRRRR=RR>hRz1hQt q75),t2
RRRRRRRRRRRRhRR 1W_QRZ =h>R 1W_Q2Z 2R;
R8CMRMVkOF0HM R)1 QZ;R

RMVkOF0HM R)1 QZR)5qt1,RQ_Z )R 1:aR17p_zmBtQ_Be a2m)
RRRR0sCkRsM1_a7ztpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)
R5RRRRR R)1 QZR)5qtRRRR>R=R1zhQ th7)5qt
2,RRRRRRRRRRRRR RhWQ_1Z= R>QR1Z) _ D1'C0MoE;22
CRRMV8Rk0MOHRFM)Q 1Z
 ;
-RR-============================================================================R

RR--QR8:7
34RkRVMHO0FaMRmh_Qa  t)qR5):tRR71a_mzpt_QBea BmR)2skC0shMRq)azqHpR#R
RLHCoMR
RRCRs0MksR_amQ hat5 )zQh1t7h 5tq)2
2;RMRC8kRVMHO0FaMRmh_Qa  t)
;
R-R-R:Q8Rd73
VRRk0MOHRFMa1F_0F8poeHOCFO0sqR5)Rt,1 QZRh:Rq)azqRp2skC0s1MRap7_mBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17m_pt_QBea Bm5)Razm_ht1Qh5 7qR)tRR=>q,)t
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR1Z= R>QR1Z2 2;R
RCRM8VOkM0MHFR_aF1p08FOoHe0COF
s;
-RR-8RQ:3R76R
RVOkM0MHFR_aF1z08pHFoOOeC0RFs5tq),QR1Z: RRahqzp)q2CRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)Razm_ht1Qh5 7qR)tRR=>q,)t
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR1Z= R>QR1Z2 2;R
RCRM8VOkM0MHFR_aF1z08pHFoOOeC0;Fs
R
RVOkM0MHFR_aF1p08FOoHe0COF5sRqR)t:qRhaqz)p1;RQ_Z )R 1:aR17m_pt_QBea Bm
)2RRRRskC0s1MRap7_mBtQ_Be aRm)HR#
RoLCHRM
RsRRCs0kMaR17m_pt_QBea Bm5)Razm_ht1QhR 75tq)R>R=Rtq),R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR1 QZRR=>1 QZ_1) 'MDCo20E2R;
R8CMRMVkOF0HMFRa_810pHFoOOeC0;Fs
R
RVOkM0MHFR_aF1z08pHFoOOeC0RFs5tq)Rh:Rq)azqRp;1 QZ_1) R1:Raz7_pQmtB _eB)am2R
RRCRs0MksR71a_mzpt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR71a_mzpt_QBea Bm5)Razm_ht1QhR 75tq)R>R=Rtq),R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRZ1Q >R=RZ1Q  _)1C'DMEo02
2;RMRC8kRVMHO0FaMRF0_18FzpoeHOCFO0s
;
CRM8b	NONRoCL$F8Rvhz B)Q_71a_1zhQ th7
;

