--$Header: //synplicity/mapgw/designware/dw01.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---a-RHC0DRRRRR:RRRj8I4E3P8-
-R#7CHRoMRRRRRB:RFNM0HRM#.L4RNO#HR#7CHWoMNRsCObFlFMMC0
#R-B-RFNlbMR$RR:RRRM1$bODHHR0$Q3MO
R--7CN0RRRRRRRR:kRqo6R.,jR.j
UR-q-RkF0EsRRRR:RRRD1CPRNl)-
-RseC#MHFRRRRRd:R3-4
--
--------------------------------------------------------------------------------------------------D

HNLssQ$R ,  7)Wq W,7j
4;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#Rq7W)7 3WObN	CNo#D3NDk;
#7CRW3j474Wj_lOFbCFMM30#N;DD
M
C0$H0R_7WMlFsR
H#oCCMsRHO5_
NI0H8ERR:uQm1a QeRR:=U#;
s_OEI8HMRu:Rma1QQRe :U=R;G
CbH_I8R0E:mRu1QQae: R=;Rc
bCG_sO0RQ:Rhta  :)R=
Rj2
;
b0FsRN5
RH:RM0R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;C_GbF#VVC:0RRRHM#_08DHFoOC_POs0F5bCG_8IH04E-RI8FMR0Fj
2;M8F_CO0C0F:Rk#0R0D8_FOoH;P
FVRD:FRk0#_08DHFoOL;
:kRF00R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;C_GbN:8[R0FkR8#0_oDFHPO_CFO0sG5CbH_I8-0E4FR8IFM0R
j22
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINC0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WMlFsRC:RM00H$#RHRC"IN;	"
C

M78RWF_Ms
l;
s
NO0EHCkO0ssCR0FDRVWR7_sMFl#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;

oLCH
M
CRM8s;0D
-

---------------------------------------------------------------------------------------------
-
DsHLNRs$Q   ,q7W)7 ,W;j4
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCWR7q3) 7NWbOo	NCN#3D
D;kR#C74Wj3j7W4F_OlMbFC#M03DND;C

M00H$WR7_sMFlM_s8#RH
MoCCOsHRN5
_8IH0:ERR1umQeaQ =R:R;4n
O#sEH_IM:8RR1umQeaQ =R:R
c;C_GbI0H8ERR:uQm1a QeRR:=cL;
_8IH0:ERR1umQeaQ =R:R;4j
bCG_sO0RQ:Rhta  :)R=
Rj2
;
b0FsRN5
_olNRH:RM0R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;b_F#F#VVC:0RRRHM#_08DHFoOC_POs0F5bCG_8IH04E-RI8FMR0Fj
2;#O0H	L$_H:0RRRHM#_08DHFoON;
_o#HMRR:H#MR0D8_FOoH;M
s8F_l8:CRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;F
b#s_CsF:Rk#0R0D8_FOoH;F
M_08CC:O0R0FkR8#0_oDFH
O;LF:Rk#0R0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R;j2
#bF:kRF00R#8F_Do_HOP0COFCs5GIb_HE80-84RF0IMF2Rj

2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsNC
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRVWR7_sMFlM_s8RR:CHM00H$R#IR"C"N	;C

M78RWF_Mssl_M
8;
ONsECH0Os0kC0RsDVRFR_7WMlFs_8sMR
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;





--------------------------------------------------------------------------------------------
--
LDHs$NsR Q  W,7q,) 74Wj;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#7CRW q)3b7WNNO	o3C#N;DD
Ck#Rj7W4W37jO4_FFlbM0CM#D3ND
;
CHM007$RW_j4#sN0MH8R#o

CsMCH5ORR8IH0:ERR1umQeaQ =R:R
U;l_#LFRk0:qRhaqz)p=R:R
n;D_#LFRk0:qRhaqz)p=R:R2.R;b

FRs05HR8MRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR20;
ORR:H#MR0D8_FOoH;N
#0RR:H#MR0D8_FOoH;M
s8RR:H#MR0D8_FOoH;P
FRF:Rk#0R0D8_FOoH;F
8k:0RR0FkR8#0_oDFHPO_CFO0s#5lLk_F0#-DLk_F0FR8IFM0R
j22
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4N_#08sMRC:RM00H$#RHRC"IN;	"
8CMRj7W4N_#08sM;N

sHOE00COkRsCsR0DF7VRW_j4#sN0MH8R#R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;C
Lo
HM
8CMRDs0;


-------------------------------------------------------------------------


DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83DSD;
M
C0$H0R_7W#VEH0RCsH
#
SCSoMHCsOS5
SNS80IN_HE80Su:Rma1QQRe :U=R;S
SRRRR#IE_HE80Su:Rma1QQRe :d=R;S
SSPHM_8lFCRS:Q hatR ):j=R
SSS2
;
SFSbsS05
SSS8NN0_SHM:MRHR8#0_oDFHPO_CFO0sN580IN_HE80-84RF0IMF2Rj;S
SS08NNO_0SH:RM0R#8F_Do;HO
SSS#SES:MRHR8#0_oDFHPO_CFO0sE5#_8IH04E-RI8FMR0Fj
2;S#SSEO_0R:RSRRHM#_08DHFoOS;
SES#_8lFCRS:H#MR0D8_FOoH;S
SS08NNk_F0F:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0FjS2
S;S2S-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7#W_E0HVC:sRR0CMHR0$H"#RI	CN"S;
SSSSSSSSSRSR
8CMR_7W#VEH0;Cs
N

sHOE00COkRsCsR0DF7VRWE_#HCV0s#RH
R

R-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM


CRM8s;0D
-

-------------------------------------------------------------------------------------------------
--
S
SSHSDLssN$CRHC
C;
SSSSCk#RCHCC03#8F_Do_HO4c4n3DND;S
SS#SkCCRHC#C30D8_FOoH_#kMHCoM8D3NDS;
SkSS#HCRC3CCMCkls_HO#308N;DD
S

SCSSM00H$WR7jO4_#HNR#S

SSSSoCCMsRHO58IH0HE:Mo0CC=s:US2;SRRR-I--HE80SRH#NCRoMHCsONRbsCNl0RCs0#FRbHCOVM$RkClLsVRFR0LH#FRVsER0CMRHb#k0R8NMR0Fkb#k0
SSSSFSbs
05SSSSSNSSSSS:SRHM#_08DHFoOC_POs0FRH5I8-0E4FR8IFM0R;j2
SSSSSSSL:SSSMSHR8#0_oDFHPO_CFO0sIR5HE80-84RF0IMF2Rj;S
SSSSSSSOS:HSSM0R#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S;
SSSSSHSOSSS:SRHM#_08DHFoOS;
SSSSSkS#l:SSSkSF00R#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S;
SSSSSNSOsSs$:FSSk#0R0D8_FOoH_OPC0RFs58IH04E-RI8FMR0Fj
2;SSSSSOSSF:SSSkSF00R#8F_Do
HO
SSSSRSS2S;
S-SS-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRSSSSRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRSSSSRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV74Wj_NO#RC:RM00H$#RHRC"IN;	"
S
SSCSSM78RW_j4O;#N
S
SSNSSsHOE00COkRsCsR0DF7VRW_j4OR#NH
#
SSSS-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRSSSR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRSRSSR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
SSSSLSSCMoH
SSSSSSS
SSSS
SSSSSSSMSC80RsDR;S
-

--------------------------------------------------------------------------------
D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
M
C0$H0Rj7W4#_NE#RH
o
SCsMCH
O5SqSS_8IH0RER:FRb#HH0P:CR=;RU
SSS1I]_HE80Rb:RF0#HHRPC:U=R
RSSR;R2
b
SF5s0RS
SSSqRSH:RM0R#8F_Do_HOP0COFqs5_8IH04E-RI8FMR0Fj
2;S7SSq_aqa:BRRRHM#_08DHFoOS;
S]S1R:SSRRHM#_08DHFoOC_POs0F5_1]I0H8ER-48MFI0jFR2S;
S]S1_RaBSH:RM0R#8F_Do;HO
SSSA:SSR0FkR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2S
S2
;
SR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jN4_#:ERR0CMHR0$H"#RI	CN"
;
CRM874Wj_EN#;


NEsOHO0C0CksRDs0RRFV74Wj_EN#R
H#
HS#oDMNR_#E.:#RR8#0_oDFHPO_CFO0s]51_8IH04E-RI8FMR0Fj
2;
RRR-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
M
C80RsD
;
---------------------------------------------------------------------------------------------


DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7_bOl_R8GHS#
oCCMs5HO
SSSI0H8ERRRRM:RNs0kN:DR=;Rc
SSSbI4_HE80RM:RNs0kN:DR=
R.S2SS;b
SF5s0RS
SSSNRSH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSSLRSH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSR0OSRS:H#MR0D8_FOoH;S
SSD8bG:RSRRHM#_08DHFoOS;
S0SD4:RSR0FkR8#0_oDFH
O;SCSSJS4R:kRF00R#8F_Do;HO
SSSoR04SF:Rk#0R0D8_FOoH;S
SS.D0RRS:FRk0#_08DHFoOS;
SJSC.:RSR0FkR8#0_oDFH
O;SoSS0S.R:kRF00R#8F_Do
HOS;S2
-
S-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7OW_l8b_GRR:CHM00H$R#IR"C"N	;C

M78RWl_ObG_8R
;
NEsOHO0C0CksRDs0RRFV7OW_l8b_GHRR#
R
R-RR-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-
----------------------------------------------------------------------------------
-
DsHLNRs$R Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DDSC

M00H$WR7j84_CHOR#o
SCsMCH
O5SISSHE80RM:RNs0kN:DR=
RcS2SS;S
Sb0Fs5SR
SRSqRRRR:MRHR0S#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S;
SzS1vRRR:kRF00R#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S
SS
2;SR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7j74_C:ORR0CMHR0$H"#RI	CN"C;
M78RW_j47;CO
s
NO0EHCkO0ssCR0FDRVWR7j74_CHOR#RR
R-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0RD;R


-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs74Wj_OHMR========================
=
DsHLNRs$R Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DDSC

M00H$WR7jH4_MHOR#o
SCsMCH
O5SISSHE80RM:RNs0kN:DR=
RcS2SS;S
Sb0Fs5SR
SRSqRRRR:MRHR0S#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S;
SzS1vRRR:kRF00R#8F_Do_HOP0COF5sRI0H8ER-48MFI0jFR2S
SS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jH4_M:ORR0CMHR0$H"#RI	CN"
;
CRM874Wj_OHM;N

sHOE00COkRsCsR0DF7VRW_j4HRMOH
#RR-RR-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;LHCoMC

Ms8R0RD;R
R
-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs74Wj_8q8R========================
=
DsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#QCR 3  #_08DHFoOM_k#MHoCN83D
D;
0CMHR0$74Wj_8N8R
H#SMoCCOsH5S
SS8IH0:ERR0MNkDsNRU:=
SSS2S;
SsbF0
5RSqSSSRR:HRMRS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSARRRRH:RMSRR#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj
2;S1SSzRvR:kRF0#RS0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SQSBR:RRRRHMR0S#8F_Do;HO
SSSBRmRRF:RkS0R#_08DHFoOS
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W48_N8RR:CHM00H$R#IR"C"N	;M
C8WR7jN4_8
8;
ONsECH0Os0kCsRR0mDRwWR7jN4_8H8R#R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsDR;R
-R
-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j4Q7hB =BR========================
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HOkHM#o8MC3DND;


CHM007$RW_j4H8MOCHOR#o
SCsMCH
O5SISSHE80RM:RNs0kN:DR=
RUS2SS;S
Sb0Fs5S
SSSqS:MRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSBQh_B7 SH:RM#RS0D8_FOoH;S
SSv1zRRS:FRk0S8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0RRj2S
SRS2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV74Wj_OHM8RCO:MRC0$H0RRH#"NIC	
";CRM874Wj_OHM8;CO
s
NO0EHCkO0ssCR0FDRVWR7jH4_MCO8O#RHRR
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoM
R
CRM8s;0D
-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7j14_z=AR========================
H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HOkHM#o8MC3DND;C

M00H$WR7j#4_kHLR#o
SCsMCH
O5SISSHE80RM:RNs0kN:DR=
RUS2SS;b
SF5s0
qSSSH:RM#RS0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S:ASRRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
BSSQRS:HSMR#_08DHFoOS;
SSBm:kRF0#RS0D8_FOoH;S
S7wQw:kRF0#RS0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2SR
S
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4k_#LRR:CHM00H$R#IR"C"N	;M
C8WR7j#4_k
L;
ONsECH0Os0kCsRR0mDRwWR7j#4_kHLR#R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;
-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs74Wj_7q71RzA=========================H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HOkHM#o8MC3DND;C

M00H$WR7jN4_8k8#L#RH
CSoMHCsOS5
SHSI8R0E:NRM0NksD=R:RSU
S;S2
FSbs
05SSSqSH:RM#RS0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SSAS:MRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SBSQS:MRHR0S#8F_Do;HO
qSS717_z:ASRRHMS8#0_oDFH
O;SmSBSRS:FRk0S8#0_oDFH
O;SzS1vRRRRRR:FRk0S8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0RRj22
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W48_N8L#kRC:RM00H$#RHRC"IN;	"
M
C8WR7jN4_8k8#L
;
qEsOHO0C0CksR0RsDwRmRj7W48_N8L#kR
H#R-RR-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCH
M
CRM8s;0D
-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7jN4_LN#PD=R======================
==
LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;
CHM007$RW_j4NPL#NHDR#C
oMHCsOS5
S8IH0:ERR0MNkDsNRR:=UR
SR2RR;F
bs
05SSqS:MRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;q
SAq1epRS:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjS2
2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4L_N#DPNRC:RM00H$#RHRC"IN;	"
M
C8WR7jN4_LN#PD
;
NEsOHO0C0CksRDs0RRFV74Wj_#NLPRNDRRH#
RRR-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCRR
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";
R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM

RRCRM8s;0D
-

-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j4O.lbR========================D=
HNLssQ$R ;  
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
M
C0$H0Rj7W4l_ObH.R#o
SCsMCH
O5SISSHE80RM:RNs0kN:DR=
RUS2SS;b
SF5s0
SSSq:SSRMRHR0S#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SSSAS:HRRM#RS0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S SpT:SSRMRHR0S#8F_Do;HO
SSSaSBS:HRRM#RS0D8_FOoH;S
SS_t t:aSRkRF0#RS0D8_FOoH;S
SS_pap: SRkRF0#RS0D8_FOoH
2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV74Wj_bOl.RR:CHM00H$R#IR"C"N	;C

M78RW_j4O.lbR
;
NEsOHO0C0CksRDs0RRFV74Wj_bOl.HRR#
R
R-RR-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsRR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"
;
-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCHCM
Ms8R0
D;
-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7jO4_lRbn=========================H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
0CMHR0$74Wj_bOln#RH
oSSCsMCH
O5SSSSI0H8ERR:MkN0sRND:U=R
SSSS
2;SFSbs50R
SSSqRS:RRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSARS:RRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSa:BSRMRHR0S#8F_Do;HO
SSSt: SRkRF0#RS0D8_FOoH;S
SSSta:FRRkS0R#_08DHFoOS;
SaSpSR:RFRk0S8#0_oDFH
O;SpSS RS:R0FkR0S#8F_Do;HO
SSSh: SRkRF0#RS0D8_FOoH;S
SSS T:FRRkS0R#_08DHFoOS
SS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jO4_lRbn:MRC0$H0RRH#"NIC	
";
8CMRj7W4l_Ob;nR
s
NO0EHCkO0ssCR0FDRVWR7jO4_lRbnRRH#
R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsDR;
RRRRR-R
-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRW_j4l_kGNRM$=========================D

HNLssQ$R ;  
Ck#R Q  a317m_pt_QB4c4n3DND;D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j4l_kGNRM$HR#
RRRRRoRRCsMCH
O5RRRRRRRRRRRRRRRRRRRRRRRRqH_I8R0ER:RRR#bFHP0HC=R:R;d.
RRRRRRRRRRRRRRRRRRRRRRRRp1 _8IH0RER:FRb#HH0P:CR=;R.
RRRRRRRRRRRRRRRRRRRRRRRRXvz_8IH0RER:FRb#HH0P:CR=
RURRRRRRRRRRRRRRRRRRRRRRRR2R;
RRRRRRRRRRRRRbRRF5s0
RRRRRRRRRRRRRRRRRRRRRRRRRqRRRRRRR:RHRMRR8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2R;
RRRRRRRRRRRRRRRRRRRRR1RR RpRR:RRRMRHR#RR0D8_FOoH_OPC05Fs1_ pI0H8ER-48MFI0jFR2R;
RRRRRRRRRRRRRRRRRRRRRvRRzRXRR:RRRkRF0#RR0D8_FOoH_OPC05Fsv_zXI0H8ER-48MFI0jFR2R
RRRRRRRRRRRRRRRRRRRRRR;R2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7jl4_kNG_M:$RR0CMHR0$H"#RI	CN"
;
CRM874Wj_Glk_$NM;


NEsOHO0C0CksRp)aRRFV74Wj_Glk_$NMR
H#
R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C8aR)p
;
-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs74Wj_O8CFR8C=========================D

HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j48FCO8HCR#SR
oCCMs5HO
SSSI0H8ERR:MkN0sRND:4=R
SSS2S;
b0Fs5S
Sq:RSRRHMS8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
ASSRRS:FRk0S8#0_oDFHPO_CFO0s*5.*8IH04E-RI8FMR0FjS2
S
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4C_8OCF8RC:RM00H$#RHRC"IN;	"
8CMRj7W4C_8OCF8;N

sHOE00COkRsCsR0DF7VRW_j48FCO8HCR#R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsDR;R
=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj7W4s_bHOCMR========================
=

H
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HON0sHED3ND
;
CHM007$RW_j4bCsHMHOR#o
SCsMCH
O5SqSS_8IH0RERR:RRR#bFHP0HC=R:R
U;SQSShX7 _8IH0:ERR#bFHP0HC=R:RSU
S;S2RS
Sb0Fs5S
SSSqRSR:RHRMRS8#0_oDFHPO_CFO0s_5qI0H8EFR8IFM0R;42RR--vHF8V8HCRRL$1PCDN0lRFNRl0ROEPHCsDRFoObFlFMMC0CR8OsDNNF0HMS
SS7Qh :XSRkRF0#RS0D8_FOoH_OPC05FsQ h7XH_I8-0E4FR8IFM0R
j2S2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV74Wj_HbsCRMO:MRC0$H0RRH#"NIC	
";
8CMRj7W4s_bHOCM;N

sHOE00COkRsCsR0DF7VRW_j4bCsHMHOR#R
RRR--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;


LHCoMC

Ms8R0
D;
=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFRj7W4H_LMOCMR========================
=
SH
DLssN$ RQ 
 ;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#R Q  03#8F_Do_HON0sHED3ND
;
CHM007$RW_j4LCHMMHOR#C
oMHCsOS5
SIq_HE80Sb:RF0#HHRPC:U=R;S
Sq)77_8IH0RER:FRb#HH0P:CR=
RcSSSS2
;RSFSbs
05SqSSSRR:RRHMR#RR0D8_FOoH_OPC05FsqH_I8-0E4FR8IFM0R;j2
SSSq)77RR:RFRk0R0R#8F_Do_HOP0COFqs57_7)I0H8ER-48MFI0jFR2S
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4H_LMOCMRC:RM00H$#RHRC"IN;	"
M
C8WR7jL4_HMMCO
;
NEsOHO0C0CksRDs0RRFV74Wj_MLHCRMOQR1
R-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs74Wj_EL#R========================D=
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM007$RW_j4LR#EH
#RSMoCCOsH5S
SSIq_HE80RRR:bHF#0CHPRR:=.S;
S]S1_8IH0:ERR#bFHP0HC=R:RS4
S;S2
bSSF5s0
SSSqRS:RRHMS8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2S;
S]S1RRR:RRHMS8#0_oDFHPO_CFO0s]51_8IH04E-RI8FMR0Fj
2;SASSSR:RFRk0S8#0_oDFHPO_CFO0s_5qI0H8ER-48MFI0jFR2S
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFRj7W4#_LERR:CHM00H$R#IR"C"N	;M
C8WR7jL4_#
E;
ONsECH0Os0kC0RsDFRRVWR7jL4_#HER#R

R-R-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;-

-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoMC

Ms8R0
D;




