-- $Header: //synplicity/mapgw/mappers/xilinx/lib/generic/gen_generic/cmp_eq.vhd#1 $
@E


DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;
0CMHR0$CCJ_DCClMH0R#R
RRFRbsN05jL,RjN,R4L,R4D,R0RHM:MRHR8#0_oDFH
O;RRRRRRRRRRRRRFD0kR0:FRk0#_08DHFoO
2;CRM8CCJ_DCClM
0;
s
NO0EHCkO0sCCRJFMRVJRC_CCDl0CMR
H#So#HMRND0:4RR8#0_oDFH
O;SO
SFFlbM0CMRXvzBpY_
SRSb0FsRR5
RSRSSRpm:kRF00R#8F_Do;HO
RRRSBSSQRR:H#MR0D8_FOoH;R
RRSSS7:QRRRHM#_08DHFoOR;
RSRSS:1RRRHM#_08DHFoOS
RS
2;S8CMRlOFbCFMM
0;SN--0H0sLCk0RNLDOL	_FFGRVzRvXRBY:FROlMbFCRM0H0#Rs;kC
oLCHSM
0<4R=MR5F50RNG4RFLsR4R22NRM850MFRj5NRsGFR2Lj2R;
RlRRkHG_MR#0:zRvX_BYpR
RRRRRRFRbsl0RN1b5RR=>0R4,
RRRRRRRRRpm=D>R00Fk,R
RRRRRRQRBRR=>DM0H,R
RRRRRRQR7RR=>'24';M
C8JRCM
;

LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
M
C0$H0R_CJClDCC_M0FLMCHH0R#R
RRFRbsN05jL,RjD,R0RHM:MRHR8#0_oDFH
O;RRRRRRRRRRRRRFD0kR0:FRk0#_08DHFoO
2;CRM8CCJ_DCClMF0_MHCL0
;

ONsECH0Os0kCJRCMVRFR_CJClDCC_M0FLMCHH0R##
SHNoMD4R0R#:R0D8_FOoH;

SSlOFbCFMMv0RzYXB_Rp
SFSbs50R
RRRSpSSmRR:FRk0#_08DHFoOR;
RSRSSRBQ:MRHR8#0_oDFH
O;RSRRSQS7RH:RM0R#8F_Do;HO
RRRS1SSRH:RM0R#8F_Do
HOR2SS;C
SMO8RFFlbM0CM;-
S-0N0skHL0LCRD	NO_GLFRRFVvBzXYRR:ObFlFMMC0#RHRk0sCL;
CMoH
4S0RR<=MRF05RNjGRFsL;j2
RRRRGlk_#HM0RR:vBzXY
_pRRRRRRRRb0FsRblN5=1R>4R0,RR
RRRRRpRRm>R=RFD0k
0,RRRRRRRRB=QR>0RDH
M,RRRRRRRR7=QR>4R''
2;CRM8C;JM



DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;
0CMHR0$B_vu HTR#R
RRCRoMHCsOH5I8R0E:MRH0CCos=R:4;d2
RRRRsbF0:5qRRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRR:RARRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRRTR RF:Rk#0R0D8_FOoH2C;
MB8Rv u_T
;

ONsECH0Os0kCCRODDD_CDPCRRFVB_vu HTR#V

k0MOHRFMVOkM_sCsFCs5JH_I8R0E:MRH0CCoss2RCs0kM0R#soHMR
H#LHCoMR
RH5VR5_CJI0H8E=R>RRU2NRM85_CJI0H8E=R<R2nc2ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5s"Cs"Fs2R;
R8CMR;HV
8CMRMVkOs_Cs;Fs
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;0
N0LsHkR0CoCCMsFN0sC_sb0FsRRFVODCD_PDCC:DRRONsECH0Os0kC#RHRMVkOs_Cs5FsI0H8E
2;
FSOMN#0MH0R0NCs0MHFRH:RMo0CC:sR=IR5HE802;/.
FSOMN#0Ms0RCHlNMs8CRH:RMo0CC:sR=IR5HE802FRl8;R.
RRRRo#HMRND8NN0_b0lR#:R0D8_FOoH_OPC0RFs58IH0-ERR84RF0IMF2Rj;R

RORRFFlbM0CMR_CJClDCCRM0HR#
RRRRRbRRF5s0NRj,LRj,NR4,LR4,DM0H:MRHR8#0_oDFH
O;RRRRRRRRRRRRRRRRRFD0k:0RR0FkR8#0_oDFH;O2
RRRR8CMRlOFbCFMM
0;
FSOlMbFCRM0CCJ_DCClMF0_MHCL0#RH
RRRRRRRRsbF0j5N,jRL,0RDHRM:H#MR0D8_FOoH;R
RRRRRRRRRRRRRRDRR00FkRF:Rk#0R0D8_FOoH2R;
RCRRMO8RFFlbM0CM;#
RHNoMD4R0R#:R0D8_FOoH;C
Lo
HMSRzj:VRH5HRI8R0E>2R4RMoCC0sNCL
SCMoH
RRRR4zjRC:RJD_CCMlC0R
RRRRRRRRRRRRRRFRbsl0RN
b5SSSSN=jR>5RqjR2,
RRRRRRRRRRRRRRRRRLj=A>R5,j2
SSSSRN4=q>R5,42RR
RRRRRRRRRRRRRR4RLRR=>A254,R
RRRRRRRRRRRRRR0RDH=MR>jR''R,
RRRRRRRRRRRRRDRR00FkRR=>8NN0_b0l52j2;C
SMo8RCsMCN;0C
R
RRRRRRSR
z:4RR5HVR8IH0=ERRR42oCCMsCN0
CSLo
HMSTS RR<=q25jRFGMs5RAj
2;S8CMRMoCC0sNC
;
RRRRz:.RRsVFR0LH_8HMCHGRMRR405FRHs0CNF0HMRR-4R2RoCCMsCN0
RRRRRRRRoLCHRM
RRRRRRRRRzRR.:4RR_CJClDCC
M0RRRRRRRRRRRRRRRRb0FsRblN5S
SSjSNRR=>q*5.L_H0HCM8GR2,
RRRRRRRRRRRRRRRRRLj=A>R5L.*HH0_MG8C2S,
SNSS4>R=R.q5*0LH_8HMC+GRR,42RR
RRRRRRRRRRRRRR4RLRR=>A*5.L_H0HCM8GRR+4
2,RRRRRRRRRRRRRRRRDM0HRR=>8NN0_b0l50LH_8HMC-GRR,42
RRRRRRRRRRRRRRRRFD0k=0R>NR800N_lLb5HH0_MG8C2
2;RRRRRRRRCRM8oCCMsCN0;S

z:dRR5HVRlsCN8HMC=sRRN4RMI8RHE80R4>R2CRoMNCs0SC
LHCoMS
SzRd4:JRC_CCDl0CM_CFML
H0SbSSFRs0l5Nb
SSSSRNj=q>R58IH0-ER4
2,SSSSL=jR>5RAI0H8ERR-4
2,SSSSDM0HR8=>N_0N05lbHs0CNF0HMRR-4
2,SSSSDk0F0>R=R204;S
SSTS RR<=M5F00;42
MSC8CRoMNCs0
C;
RRRRRRRRz
ScRR:HsV5CHlNMs8CRj=RR8NMR8IH0RER>2R4RMoCC0sNCL
SCMoH
RRRRTS RR<=M5F08NN0_b0l5CH0sHN0F-MRR242;
R
S8CMRMoCC0sNC
;
CRM8RDOCDC_DP;CD








