@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)]a_q1h7] qi"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
`8HVCmVReqp_1)1 ah_m
R
RsRCoV#Hs0C_sJ
;
RDRNI#N$RR@@5#bFCC8oR	OD2CRLo
HMRRRRH5VR`pme_1)  1a_Qqthp=R!RL4'jL2RCMoH
RRRRHRRVV55H0s#_JsCRV^RH0s#_JsC2=R=RL4'jL2RCMoH
RRRRRRRRRHV5JsC2R
RRRRRRRRRV#Hs0C_sJ=R<RL4'4R;
RRRRRCRRMR8
RRRRRCRRDR#CLHCoMR
RRRRRRRRRV#Hs0C_sJ=R<RL4'jR;
RRRRRCRRMR8
RRRRR8CM
RRRR#CDCR
RRRRRV#Hs0C_sJ=R<RL4'jR;
R8CM
R
RbbsFC$s0R1q1 _)a]7qh1i]q B_qiQ_vhY_BB_p uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RFfs#sC5CRJ2|R->5f!5sCF#5	NO2R22rH*lMO_N	$_OO9DC;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)]a_q1h7] qi_iqB_Xvq_BBYpu _;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
Rf#sFCC5sJ&2R&!R5f#sFCO5N	R22|R->
5RRy4yr:N5lGO_N	$_OORDC>RRj?NRlGO_N	$_OORDC:2R.9fR5sCF#5	NO2|R|Rs5fF5#Cs2CJRR&&5JsC_F8sb=R=RL4'42222R;
R8CMbbsFC$s0

RRRsRbFsbC0q$R1)1 aq_]h]71q_i q_Biv_qXpt hau]_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
Rf#sFCO5N	|2R-5>RN2O	r:*45GlN_	NO_MDCoR0E>RRj?NRlGO_N	C_DMEo0R.:R2RR9yRy45O!N	
2;RMRC8Fbsb0Cs$
R
RsRbFsbC0q$R1)1 aq_]h]71q_i )_ T7u)m_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RsRfF5#Cs2CJR>|-RC5sJ4r*:2f9RjyyRFfs#NC5O;	2
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 aq_]h]71q_i vazpQ up_T) _
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RFRM05R5f#sFCC5sJ&2R&NR!OR	2yRy45JsCRR&&!	NO2*Rrj9:fRR
RyRy45C!sJ&R&RO!N	r2R*f4:9yRy4fR5sCF#5JsC2;22
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 aq_]h]71q_i )_ T71 q1a )_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RfR5sCF#5	NO2&R&RC5sJR22|R->5ryyjC:8NC##sO0_F0kM9s5!C2J2;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)]a_q1h7] qi_iqB_aWQ]amz_T) _)wQ1)a_ uT_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
Rf#sFCO5N	|2R-5>RV#Hs0C_sJ|R|RJsC2R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)a]7qh1i]q B_qiQ_Waz]ma _)Tz_1AT1 za h_T) _
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RVRfC5DDN2O	R>|-RFfs#sC5CRJ2IEH0H5MR!	NORjr*:Rf9yRy4N2O	;R
RCbM8sCFbs
0$
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRsRbFsbC0q$R1)1 aq_]h]71q_i )_ TXuZ_;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRfR!HM#k	IMFMs5RC2JR;R
RRMRC8Fbsb0Cs$R

RbRRsCFbsR0$q 11)]a_q1h7] qi_iqB__XZuR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R!RRfkH#MF	MIRM5NRO	2R;
RCRRMs8bFsbC0R$
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRHRRVlR5HNM_OO	_$CODRj>R2CRLoRHM:_RNNC##sE0_N#M8ECN	_	NO_MlH_OO$DRC
RRRRRRRRRqq_1)1 aq_]h]71q_i q_Biv_QhBpYB :_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)]a_q1h7] qi_iqB_hvQ_BBYpu _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5O"q	IMFDoC8C#RN#0CsCL8RCsVFCDRCNCb#RRFV#ObCHCVH8HRlMkHllHRlMO_N	$_OORDCOD$OCV#RsRFlskCJC"#02R;
RRRRRCRRMR8
RRRRRHRRVlR5NNG_OO	_$CODRj>R2CRLoRHM:_RNNC##sE0_N#M8ECN	_	NO_GlN_OO$DRC
RRRRRRRRRqq_1)1 aq_]h]71q_i q_Biv_qXBpYB :_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)]a_q1h7] qi_iqB_Xvq_BBYpu _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5O"q	IMFDoC8C#RHR0MFR#N#CCs08HRI0MEHRC#bOHHVCl8RNlGHkllRNNG_OO	_$CODROO$DRC#VlsFRJsCk0C#"
2;RRRRRRRRC
M8RRRRRRRRH5VR5GlN_	NO_MDCoR0E>4=R2L2RCMoHRN:R_#N#C_s0E8NM#	ENCO_N	N_lGC_DMEo0
RRRRRRRRqRR_1q1 _)a]7qh1i]q B_qiq_vX _ph]ta_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_]h]71q_i q_Biv_qXpt hau]_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5k"7sHN0FFMRVFROMM0Hk#FkR#N#CCs080R#NR0CFNVROF	MI8DCoPCRHNFD0RC##ObCHCVH8NRlGkHllORN	N_lGC_DMEo0ROO$D"C#2R;
RRRRRCRRMR8
RRRRRHRRV8R5C#N#C_s0OMFk0RR>jL2RCMoHRN:R_#N#C_s0E8NM#	ENCC_sJC_8NC##sR0
RRRRRRRRRqq_1)1 aq_]h]71q_i )_ T71 q1a )_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_]h]71q_i )_ T71 q1a )_
u2RRRRRRRRRDRC#FCRPCD_sssF_"057Nks0MHFRRFVO0FMHFMkkN#R#s#C0RC8#00NCVRFRJsCk0C#RFPHDCN0#bR#CVOHHRC88#CN#0Cs_kOFMO0R$COD#;"2
RRRRRRRR8CM
RRRRRRRRRHV5JsC_F8sbRR>jL2RCMoHRN:R_#N#C_s0E8NM#	ENCC_sJs_8FRb
RRRRRRRRRqq_1)1 aq_]h]71q_i )_ T7u)m_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_]h]71q_i )_ T7u)m_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05)kCJCR#0H8#RC#N#CCs08CRLVCFsR	NOMDFICC8ol0CMRsNsH#PC"
2;RRRRRRRRC
M8RRRRRRRRq1_q1a )_h]q7q1]iv _zQpau_p )_ TuR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)]a_q1h7] qi_pvzapQu  _)T2_u
RRRRRRRR#CDCPRFDs_Cs_Fs0h5"CsIRCCJk#N0RsPsHCL#RCsVFCsRbCFPHks#RCCJk#H0R#ORN	IMFDoC8C28";R
RRRRRR_Rqq 11)]a_q1h7] qi_iqB_aWQ]amz_T) _)wQ1)a_ uT_:R
RRRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_]h]71q_i q_BiW]Qam_za)_ Tw1Q)a _)T2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"	qOMDFICC8oRsNsH#PCR0IHE0FkRbNRCHM8MsoRCCJk#20";R
RRRRRR_Rqq 11)]a_q1h7] qi_iqB_aWQ]amz_T) _A1z1z T _ha)_ TuR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)]a_q1h7] qi_iqB_aWQ]amz_T) _A1z1z T _ha)_ TuR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0q5"OF	MI8DCoNCRsPsHCI#RHF0EkN0RRMbC8oHMRJsCk0C#"
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR/R/GR/xOOEC	oHMRsVFRJsCRo#HM
ND
RRRRRRRRqq_1)1 aq_]h]71q_i )_ TXuZ_:R
RRRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_]h]71q_i )_ TXuZ_2R
RRRRRRDRC#FCRPCD_sssF_"05sRCJO0FMN#HMRFXRs"RZ2
;
RRRRRRRR///GxEROCHO	MVoRFNsRO#	RHNoMDR

RRRRRqRR_1q1 _)a]7qh1i]q B_qiZ_X_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)a]7qh1i]q B_qiZ_X_
u2RRRRRRRRCCD#RDFP_sCsF0s_5O"N	FROMH0NMX#RRRFsZ;"2
R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRH5VRl_HMN_O	OD$OCRR>jL2RCMoHRl:R_#N#C_s0E8NM#	ENCO_N	H_lM$_OO
DCRRRRRRRRR_Rvq 11)]a_q1h7] qi_iqB_hvQ_BBYpu _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)a]7qh1i]q B_qiQ_vhY_BB_p u
2;RRRRRRRRC
M8RRRRRRRRH5VRl_NGN_O	OD$OCRR>jL2RCMoHRl:R_#N#C_s0E8NM#	ENCO_N	N_lG$_OO
DCRRRRRRRRR_Rvq 11)]a_q1h7] qi_iqB_Xvq_BBYpu _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)a]7qh1i]q B_qiq_vXY_BB_p u
2;RRRRRRRRC
M8RRRRRRRRH5VR5GlN_	NO_MDCoR0E>4=R2L2RCMoHRl:R_#N#C_s0E8NM#	ENCO_N	N_lGC_DMEo0
RRRRRRRRvRR_1q1 _)a]7qh1i]q B_qiq_vX _ph]ta_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 aq_]h]71q_i q_Biv_qXpt hau]_2R;
RRRRRCRRMR8
RRRRRHRRV8R5C#N#C_s0OMFk0RR>jL2RCMoHRl:R_#N#C_s0E8NM#	ENCC_sJC_8NC##sR0
RRRRRRRRRqv_1)1 aq_]h]71q_i )_ T71 q1a )_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 aq_]h]71q_i )_ T71 q1a )_;u2
RRRRRRRR8CM
RRRRRRRRRHV5JsC_F8sbRR>jL2RCMoHRl:R_#N#C_s0E8NM#	ENCC_sJs_8Fbb_
RRRRRRRRvRR_1q1 _)a]7qh1i]q  _)T)_7muu_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)a]7qh1i]q  _)T)_7muu_2R;
RRRRRCRRMR8
RRRRRvRR_1q1 _)a]7qh1i]q z_vpuaQp) _ uT_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 aq_]h]71q_i vazpQ up_T) _;u2
RRRRRRRRqv_1)1 aq_]h]71q_i q_BiW]Qam_za)_ Tw1Q)a _)T:_u
RRRRRRRR#N#kRlCbbsFC$s0R15q1a )_h]q7q1]iq _BWi_Qma]z)a_ wT_Qa)1_T) _;u2
RRRRRRRRqv_1)1 aq_]h]71q_i q_BiW]Qam_za)_ T11zA  Tzh)a_ uT_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 aq_]h]71q_i q_BiW]Qam_za)_ T11zA  Tzh)a_ uT_2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRG///OxRE	COHRMoVRFssRCJ#MHoN
D
RRRRRRRRv1_q1a )_h]q7q1]i) _ XT_Z:_u
RRRRRRRR#N#kRlCbbsFC$s0R15q1a )_h]q7q1]i) _ XT_Z2_u;R

RRRRR/RR/xG/RCOEOM	HoFRVsORN	HR#oDMN
R
RRRRRR_Rvq 11)]a_q1h7] qi_iqB__XZuR:
RRRRRNRR#l#kCsRbFsbC05$Rq 11)]a_q1h7] qi_iqB__XZu
2;
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
RCRoMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RRRROCFPsC_sJ#_N#0CsC
8:RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R`55m_ep)  1aQ_1tphqRR!=4j'L2&R&RFfs#sC5C2J22R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05s_CJNC##s80CRPOFC8sC"
2;
RRRRFROP_CsN_O	NC##s80C:R
RRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52R5e`mp _)1_ a1hQtq!pR='R4LRj2&f&RsCF#5	NO2
22RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5O"N	#_N#0CsCO8RFsPCC28";R
RRMRC8R
RR8CM
R
RCoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
