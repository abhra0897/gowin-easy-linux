`ifndef ATCMSTMUX100_CONFIG_VH
`define ATCMSTMUX100_CONFIG_VH

	`define ATCMSTMUX100_ADDR_WIDTH 32
	`define ATCMSTMUX100_DATA_WIDTH 32

	`define ATCMSTMUX100_MST0_SUPPORT
	`define ATCMSTMUX100_MST1_SUPPORT
	`define ATCMSTMUX100_MST2_SUPPORT
	`define ATCMSTMUX100_MST3_SUPPORT
	`define ATCMSTMUX100_MST4_SUPPORT
	`define ATCMSTMUX100_MST5_SUPPORT
	`define ATCMSTMUX100_MST6_SUPPORT
	`define ATCMSTMUX100_MST7_SUPPORT
`endif //ATCMSTMUX100_CONFIG_VH
