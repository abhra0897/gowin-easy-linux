@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)ah  e)
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
R`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MCRCR`MV8H
H
`VV8CRpme_1q1 _)am
h
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRFbsb0Cs$1Rq1a )_eh  X)_Z;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR55!fkH#MF	MI0M5C_#0CsGb2;22
RRRR8CMbbsFC$s0
`RRCHM8V/R/Rpme_uQvpQQBaB_X]i B_wmw
M`C8RHV/m/ReXp_BB] iw_mwR

RFbsb0Cs$1Rq1a )_eh  u)_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R!H5f#	kMMMFI5#0C0G_Cb2s2R>|-RC50#C0_GRbs!4=R'2L4;R
RCbM8sCFbs
0$
oRRCsMCN
0C
RRRR#ONCbR5sCFbs_0$0C$b2R
RRRRR`pme_1q1 R)a:CRLoRHM:PRFD#_N#0Cs
RRRRRRRRqq_1)1 a _he_ )uR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)ha_ )e _
u2RRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHR0MFRpwq12 ";`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRq1_q1a )_eh  X)_Z:_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_eh  X)_Z2_u
RRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 a _he_ )uR:RR#RN#CklRFbsb0Cs$qR51)1 a _he_ )u
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rvq 11)ha_ )e __XZuN:R#l#kCsRbFsbC05$Rq 11)ha_ )e __XZu
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
