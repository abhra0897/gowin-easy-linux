--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lbj6j#/L0lbNbC/s#GHHDMDG/HoL/CPM_HCs0Gk/lDP03E48yR-f
-


---
--
-RkRvDb0HDsHCR0IHEHRbbkCLV5#RHOMRNR#CFbVRHDbCHMMHo-2
-NRas0oCRe:RHCs0G-
-
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;D

HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;C

M00H$HRwsu#0skF8OR0#HS#
oCCMs5HO
ISSHE80qRR:HCM0o;Cs
ISSHE80ARR:HCM0o
CsS
2;SsbF0
R5SRSqRH:RM#RR0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;SRSARH:RM#RR0D8_FOoH_OPC05FsI0H8E4A-RI8FMR0Fj
2;SASqRF:Rk#0R0D8_FOoH_OPC05FsI0H8EIA*HE80qR-48MFI0jFR2S
S-A-RRq*R
;S2
8CMRswH#s0uFO8k0
#;
ONsECH0Os0kCsRNORE4FwVRH0s#u8sFk#O0R
H#
RRR#MHoNNDR_GNkR#:R0D8_FOoH_OPC05FsI0H8E4q-RI8FMR0Fj
2;R#RRHNoMD_RLNRkG:0R#8F_Do_HOP0COFIs5HE80AR-48MFI0jFR2L;
CMoH
FSVs8NMqV:RFHsRNMRHR0jRFHRI8q0E-o4RCsMCN
0CSRRRVNFsM:8ARsVFRRHLHjMRRR0FI0H8E4A-RMoCC0sNCS
SqIA5HE80AN*HRH+RL<2R=5RNHRN2NRM8LL5H2S;
RCRRMo8RCsMCNR0CVNFsM;8A
MSC8CRoMNCs0VCRFMsN8
q;CRM8NEsO4
;

LDHs$NsR Q  D;
HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;#
kC RQ 1 3ap7_mBtQ_n44cD3NDb;
NNO	oeCRBumvmhh aH1R#F
OlMbFCRM0u QuA
zwSsbF0
R5SRSm:kRF00R#8F_Do;HO
QSSRH:RM0R#8F_Do
HOS
2;CRM8ObFlFMMC0
;
Ns00H0LkC$R#MD_LN_O	LRFGFuVRQAu z:wRRlOFbCFMMH0R#sR0k
C;-C-RMF8RVHRbbkCLV-

-MR 8NRLON	IsO8RFNlb0HHLD$H0RlOFbCFMM
0#CRM8evBmu mhh;a1
D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
Ck#RFPOlMbFC#M03DND;C

M00H$8RN8osCR
H#SMoCCOsH5S
SI0H8ERR:HCM0o;Cs
sSSCRoRRH:RMo0CC-sR-NRhlFCRVER0CCRDP
CDS
2;SsbF0
R5SRSqRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SRARRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SsRC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
;S2
0SN0LsHkR0C\N3sMR	\:MRH0CCosS;
Ns00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MN8R8C8so
;
NEsOHO0C0CksRONsEF4RV8RN8osCR
H#R#RRHNoMDCRs#0kDR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2L;
CMoH
RRRskC#D<0R=RRq+;RA
RRRVDFsF.Fb:FRVsRRHHjMRRR0FI0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#s;Co
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RRRRoLCHSM
s#Co:HRbbkCLVb
SFRs0l5Nb
RSRR=QR>CRs#0kD5,H2
RSRR=mR>CRs#25H
;S2
RRRCRM8oCCMsCN0RsVFDbFF.C;
MN8Rs4OE;D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3ND
;
kR#CPlOFbCFMM30#N;DD
M
C0$H0RFVDFHsR#R
RRRRRRRRRRRRRRCRoMHCsO
R5SISSHE80QRhR:MRH0CCos=R:R;gj
SSSI0H8EamzRH:RMo0CC:sR=cR6;S
SSlMkLRCsRRR:HCM0oRCs:6=R;S
SS8HMCRGRR:RRR0HMCsoCR4:=
RRRRRRRRRRRRRRRR
2;RRRRRRRRRRRRRRRRb0FsRR5
RRRRRRRRRRRRRRRRRQRRM0bkRRR:RRHM#_08DHFoOC_POs0F58IH0hEQ-84RF0IMF2Rj;R
RRRRRRRRRRRRRRRRRRkRm00bkRF:Rk#0R0D8_FOoH_OPC05FsI0H8Eamz-84RF0IMF2Rj
RRRRRRRRRRRRRRRR
2;S0N0skHL0\CR3MsN	:\RR0HMCsoC;N
S0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C8DRVF;Fs
s
NO0EHCkO0sNCRs4OERRFVVFDFs#RHRR
RRFROlMbFCRM0Ns88CSo
RCRoMHCsO
R5SSRRS8IH0:ERR0HMCsoC;S
SSosCR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPDR
SR
2;SbRRFRs05S
SqRRR:MRHR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;S
SARRR:MRHR8#0_oDFHPO_CFO0sI5RHE80-84RF0IMF2Rj;S
SsRC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
RSR2R;
RMRC8FROlMbFC;M0
V
Sk0MOHRFM#VEH0sxCFM5H8RCG:MRH0CCoss2RCs0kMMRH0CCos#RH
RSRRsPNHDNLC0R#C:bRR0HMCsoC;L
SCMoH
RSRRC#0b=R:R
4;SRRRVRFsHMRHR04RFMRH8-CG4FRDFSb
SC#0b=R:RC#0bRR*.S;
RCRRMD8RF;Fb
RSRR0sCkRsM#b0C;R
RRMSC8ER#HxV0C;sF
O
SF0M#NRM0#VEH08N8C:sRR0HMCsoCRR:=#VEH0sxCFM5H82CG;O
SF0M#NRM0DoCME:0RR0HMCsoCRR:=I0H8E/QMMLklC
s;LHCoMV
SFFsDF4b_:FRVsRR[H4MRRR0FMLklC.s/RMoCC0sNCL
SCMoH
RSRRosC#Rq:Ns88CSo
RoRRCsMCHlORN5bR
ISSHE80RR=>DoCME#0-E0HVNC88sS,
SosCR=RR>MRH8
CGSRRR2R
SRFRbsl0RN
b5SRRRRqRRRR=>QkMb0C5DM0oE**5.[2-4-84RF0IMFCRDM0oE*5.*[2-4+H#EV80N82Cs,R
SRRRRR=AR>MRQb5k0DoCME.0**4[-RI8FMR0FDoCME50*.-*[4#2+E0HVNC88s
2,SRRRRsRRC=#R>kRm00bk5MDCo*E0[R-48MFI0DFRCEMo0[*5-+42#VEH08N8C
s2SRRR2S;
RVRRFFsDF.b_:FRVsRR	HjMRRR0F#VEH08N8C4s-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#RR:DCNLD#RHR8HMC
G;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;SRRRLHCoMR
SRRRR-m-Rkk0b0C5DM0oE*-5[4#2+E0HVNC88sR-48MFI0DFRCEMo0[*5-242RR<=
-S-RSSSSMSQb5k0DoCME.0**-5[4#2+E0HVNC88sR-48MFI0DFRCEMo0**.54[-2
2;SRRRRsRRC:o#RbbHCVLk
RSRRRRRb0FsRblN5R
SRRRRRRRRQ>R=RbQMkD05CEMo0**.54[-22+	,R
SRRRRRRRRm>R=R0mkb5k0DoCME50*[2-4+
	2SRRRR2RR;R
SRMRC8CRoMNCs0VCRFFsDF.b_;C
SMo8RCsMCNR0CVDFsF_Fb4S;
H#V_FNk#:VRHRk5MlsLCR8lFR=.RRR42oCCMsCN0
CSLo
HMSRRR-F-VsFDFb:_dRsVFRHHRMRR40DFRCEMo0E-#HNV08s8CRMoCC0sNCR
SRFRVsFDFb:_dRsVFRHHRMRR40DFRCEMo0CRoMNCs0SC
S0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RSRRoLCHSM
RRRRRCRsoR#:bCHbL
kVSRRRRbRRFRs0l5Nb
RSRRRRRRQRRRR=>QkMb0H5I8Q0Eh2-H,R
SRRRRRRRRm>R=R0mkb5k0I0H8Eamz-
H2SRRRR2RR;R
SRMRC8CRoMNCs0VCRFFsDFdb_;R
SR-R-R0mkb5k0I0H8Eamz-H#EV80N8-Cs4FR8IFM0R8IH0zEmaC-DM0oE2SR
-S-RS=S<RbQMkI05HE80Q#h-E0HVNC88sR-48MFI0IFRHE80QDh-CEMo0
2;S8CMRMoCC0sNCVRH_k#F#
N;CRM8NEsO4
;
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00N$R8s8CaCsCR
H#SMoCCOsH5S
SI0H8E:qRR0HMCsoC;S
SI0H8E:ARR0HMCsoC
;S2
FSbs50R
qSSA:RRRRHM#_08DHFoOC_POs0F58IH0*EAI0H8E4q-RI8FMR0Fj
2;SsSbFO8k0RR:FRk0#_08DHFoOC_POs0F58IH0+EAI0H8E4q-RI8FMR0FjS2
SR--ARR*q2
S;M
C88RN8aCss;CC
NR
sHOE00COkRsCNEsO4VRFR8N8CssaCHCR#R
RRMOF#M0N0ER0CoEHERR:#_08DHFoOC_POs0F5R468MFI0jFR2=R:RhBmea_17m_pt_QBea BmI)5HE80q,-4R24n;R
RRlOFbCFMMV0RDsFF
RRRRoRRCsMCH5OR
SSSI0H8ERQhRH:RMo0CC;sR
SSSI0H8EamzRH:RMo0CC;sR
SSSMLklCRsRRH:RMo0CC;sR
SSSHCM8GRRRRRR:HCM0o
CsRRRRR;R2
RRRRRRRb0FsRR5
RRRRRRRRRRRRRbQMkR0R:MRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2R;
RRRRRRRRRRRRR0mkbRk0:kRF00R#8F_Do_HOP0COFIs5HE80m-za4FR8IFM0R
j2RRRRR2RR;R
RR8CMRlOFbCFMM
0;
RRRVOkM0MHFRb8C0HEW8R0EskC0sHMRMo0CCHsR#R
RRoLCHRM
RRRRVRFsHMRHRR468MFI0jFRRFDFbH
SV0R5EHCEoHE52RR='24'RC0EMR
SRCRs0MksR4H+;C
SMH8RVR;
RRRRCRM8DbFF;R
RRsRRCs0kM;Rj
RRRCRM880CbE8WH0
E;
RRRO#FM00NMRb8C0:ERR0HMCsoCRR:=80CbE8WH0
E;RORRF0M#NRM0I0H8E:0RR0HMCsoCRR:=I0H8EIA+HE80q;+4
RRR0C$bRlDH##RHRsNsN5$R80CbER+48MFI0jFR2VRFR0HMCsoC;

RRVRRk0MOHRFMOONDhLklCRs#skC0sDMRHRl#HR#
RRRRRsPNHDNLCER0Ck_MlsLC#RR:D#Hl;R
RRoLCHRM
RRRRRC0E_lMkL#Cs5Rj2:I=RHE80qR;
RRRRRsVFRHHRMRR408FRCEb0+D4RF
FbRRRRRRRRRC0E_lMkL#Cs5RH2:0=REMC_kClLsH#5-/42.RR+5C0E_lMkL#Cs54H-2FRl82R.;R
RRRRRCRM8DbFF;R
RRRRRskC0s0MREMC_kClLs
#;RRRRCRM8OONDhLklC;s#
RR
RFROMN#0MM0RkClLs:#RRlDH#=R:RDONOlhkL#Cs;

RRVRRk0MOHRFMOONDpRHlskC0sDMRHRl#HR#
RRRRRsPNHDNLCER0CH_Dl:#RRlDH#R;
RRRRRsPNHDNLCkRMl:LRR0HMCsoC;R
RRoLCHRM
RRRRRC0E_lDH#25jRR:=jR;
RRRRRlMkL=R:R8IH0;Eq
RRRRVRRFHsRRRHM4FR0Rb8C04E+RFDFbS
R0_ECD#Hl5RH2:0=REDC_H5l#H2-4RM+Rk*lLI0H8E
0;RkSMl:LR=kRMl.L/R5+RMLklR8lFR;.2
RRRRCRRMD8RF;Fb
RRRRsRRCs0kMER0CH_Dl
#;RRRRCRM8OONDp;Hl
RR
RFROMN#0MP0RCHODlRR:D#HlRR:=OONDp;Hl
RRR#MHoNLDRHso0C:CRR8#0_oDFHPO_CFO0sC5POlDH5b8C04E+2R-48MFI0jFR2
;
LHCoMSR
L0Hos5CCI0H8E40-RI8FMR0Fj<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E4q+2S
SSSRRS&SSR5qAI0H8E4A-RI8FMR0Fj
2;RVRRFMsN8Rq:VRFsHHNRMRR40IFRHE80qR-4oCCMsCN0
LSSHso0C5C5H4N+2H*I800E-84RF0IMFNRH*8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,HRI8q0E-+HN4S2
SRSRSSSS&ARq58IH0*EA5+HN442-RI8FMR0FI0H8EHA*NS2
SRSRSSSS&mRBh1e_ap7_mBtQ_Be a5m)jH,RN
2;RCRRMo8RCsMCNR0CVNFsM;8q
R
RRsVFDbFF.F:VsRR[H4MRRR0F80CbECRoMNCs0SC
lR4:RFVDFSs
SMoCCOsHRblNRS5
SHSI8Q0Eh=RR>CRPOlDH5R[2-CRPOlDH54[-2S,
SHSI8m0Ez=aR>CRPOlDH54[+2RR-PDCOH[l52S,
SkSMlsLCR=RR>kRMlsLC#-5[4
2,SHSSMG8CRRRR=[>R
SSS2S
Sb0FsRblNRS5
SRSRQkMb0RRRRR=>L0Hos5CCPDCOH[l52R-48MFI0PFRCHODl-5[4,22
SSSRkRm00bkR=RR>HRLoC0sCC5POlDH54[+2R-48MFI0PFRCHODl25[2S
SS
2;RCRRMR8RoCCMsCN0RsVFDbFF.
;
RbRRskF8O<0R=HRLoC0sCC5POlDH5b8C04E+2R-.8MFI0PFRCHODlC58b20E2
;R
8CMRONsE
4;
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
#
kCORPFFlbM0CM#D3ND
;
CHM00v$RzRpaHS#
oCCMs5HO
NSSI0H8ERR:HCM0oRCs:g=R;S
SL8IH0:ERR0HMCsoCRR:=gS;
S8IH0RER:MRH0CCos=R:R
4US
2;SsbF0
R5SRSqR:RRRRHMR8#0_oDFHPO_CFO0sI5NHE80-84RF0IMF2Rj;S
SARRRRH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;S)Sum:7RR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R
j2S-S-R*ARRSq
2S;
Ns00H0LkC3R\s	NM\RR:HCM0o;Cs
0SN0LsHkR0C\C3slCFP__MFIMNs\RR:HCM0o;Cs
8CMRpvza
;
NEsOHO0C0CksRONsEF4RVzRvpHaR#R

RkRVMHO0F#MRkIb5HE80NI,RHE80LRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRVRHRH5I8N0ERI>RHE80L02RE
CMSCRs0MksR8IH0;EN
RRRRCRRD
#CRsSRCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRM#8Rk
b;
RRRVOkM0MHFRVHM58IH0,ENR8IH0REL:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRH5VRI0H8E<NRR8IH02ELRC0EMR
SskC0sIMRHE80NR;
RRRRR#CDCs
SCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRMH8RM
V;
RRRO#FM00NMR8IH0REq:MRH0CCos=R:RVHM5HNI8,0ERHLI820E;R
RRMOF#M0N0HRI8A0ERH:RMo0CC:sR=kR#bI5NHE80,IRLHE802
;
RORRFFlbM0CMRswH#s0uFO8k0S#
oCCMs5HO
ISSHE80qRR:HCM0o;Cs
ISSHE80ARR:HCM0o
CsS
2;SsbF0
R5SRSqRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;SRSARH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;SASqRF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2S
S-A-RRq*R
;S2
RRRCRM8ObFlFMMC0
;
RORRFFlbM0CMR8N8CssaCSC
oCCMs5HO
ISSHE80qRR:HCM0o;Cs
ISSHE80ARR:HCM0o
CsS
2;SsbF0
R5SASqRRR:H#MR0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2S;
SFbs80kORF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE+I0H8ER-48MFI0jFR2S
S-A-RRq*R
;S2
RRRCRM8ObFlFMMC0
;
R#RRHNoMD_RNNRkG:0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2R;
RHR#oDMNRNL_k:GRR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;R
RRo#HMRNDNRLRRRR:#_08DHFoOC_POs0F5HNI8*0EL8IH04E-RI8FMR0Fj
2;R#RRHNoMDCRs#0kD:0R#8F_Do_HOP0COFNs5I0H8EI+LHE80-84RF0IMF2Rj;C
LoRHM
RRR-1-RIRNbqMRN8RRAHMVRC#OC#$Ns
RRRHDVqNCsosRA:H5VRN8IH0>ERRHLI820ERMoCC0sNCR
RRRRRVDFsF.Fb:FRVsRRHHjMRRR0FL8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;S
SNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;R
RRRRRLHCoMR
SRCRso:#qRbbHCVLk
RSRRsbF0NRlbS5
RRRRRRRQ=A>R5,H2
RSRRRRRm>R=RNN_kHG52R
SR;R2
RSRRosC#RA:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RqH
2,SRRRRmRRRR=>Lk_NG25H
RSRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;b.
RRRRVRRFFsDF:b4RsVFRHHRMIRLHE80RR0FN8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:ARRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#A:NRDLRCDH4#R;R
RRRRRLHCoMR
SRCRso:#ARbbHCVLk
RSRRsbF0NRlbS5
RRRRRRRQ=q>R5,H2
RSRRRRRm>R=RNL_kHG52R
SR;R2
RRRRCRRMo8RCsMCNR0CVDFsF4Fb;R
RR8CMRMoCC0sNCVRHqsDNoACs;R

RVRHqN#lDsDCAH:RVNR5I0H8E=R<RHLI820ERMoCC0sNCR
RRRRRVDFsFNFb:FRVsRRHHjMRRR0FN8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:BRRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#B:NRDLRCDH4#R;S
SNs00H0LkC3R\s	NM\VRFRosC#:1RRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#1:NRDLRCDH4#R;R
RRRRRLHCoMR
SRCRso:#BRbbHCVLk
RSRRsbF0NRlbS5
RRRRRRRQ=q>R5,H2
RSRRRRRm>R=RNN_kHG52R
SR;R2
RSRRosC#R1:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RAH
2,SRRRRmRRRR=>Lk_NG25H
RSRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bN
RRRRVRRFFsDF:bLRsVFRHHRMIRNHE80RR0FL8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:7RRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#7:NRDLRCDH4#R;R
RRRRRLHCoMR
SRCRso:#7RbbHCVLk
RSRRsbF0NRlbS5
RRRRRRRQ=A>R5,H2
RSRRRRRm>R=RNL_kHG52R
SR;R2
RRRRCRRMo8RCsMCNR0CVDFsFLFb;R
RR8CMRMoCC0sNCVRHqN#lDsDCA
;
RwRRH0s#1b0C:HRwsu#0skF8O
0#SMoCCOsHRblNRS5
S8IH0REq=I>RHE80qS,
S8IH0REA=I>RHE80A2
S
FSbsl0RN5bR
qSSRR=>Nk_NGS,
S=AR>_RLN,kG
qSSA>R=R
NLS
2;
RRRqC88sCasC:.RR8N8CssaCSC
oCCMsRHOlRNb5S
SI0H8E=qR>HRI8q0E,S
SI0H8E=AR>HRI8A0E

S2SsbF0NRlb
R5SASqRR=>N
L,SsSbFO8k0>R=R#sCk
D0S
2;
RRRRmu)7=R<R#sCk5D0I0H8ER-48MFI0jFR2C;
MN8Rs4OE;



