--
@ER--a#EHRDVHC#RHRHIs0M0CRRHMNCMRGM0C8RC8ep]7RN0E0NRlbV#Rk0MOH#FM
R--FFM0RHLkDM0H#FRVs$R1MHbDVR$3RCaERlMkCOsHRN#0Ms8N8HR#lNkD0MHFR-
-RObN	CNoR8NMRObN	CNo
R--L$F8RRH#NHPNDDNLCMRFRsNRFD$N0L$RN##HRFVslCRHC
C3---
--R--------------------------------------------------------------------------
-----
-FRBbH$soRE0�gR4gL(R$ RQ R 3qRDDsEHo0s#RCs#CP3C8

---a-RERH##sFkOVCRHRDCHN#RM#RC#0CMHRNDb0NsRRFVQ   R810R(4jn-3d4(gg,-
-R Q  0R1NNM8se8R]R7p10$MEHC##NRuOo	NCR#3a#EHRk#FsROCVCHDR$lNR0MFR
LC-O-RFCbH8#,RF,D8RRFsHDMOk88CR0IHEFR#VN0Is0CRERN0H##RFRD8IEH0FRk0I0sH0RCM
R--blCsHH##FVMRsRFl0RECQ   RN10Ms8N87#RCsbN0MlC0a3RERH##sFkOVCRHRDCl
N$-L-RC#RkC08RFlRHblDCCRM00#EHRN#0Ms8N8MRN8NRl$CRLR#8H0LsHk80CRRHMObFlH8DC
R--VlFsRRHMNRM$lMNMC#sRFFRDMNoR#ER0CFROlDbHCV8RFRsl8#FCR0MFRDNDF8IRHOsC0-
-RO8CFHlbDHN0FFMRVER0CsRFHMoHN#DRFOksCHRVDRC3a#EHRk#FsROCVCHDR$lNRRLC
R--OHFbCV8RFHsRMP8HHN8kD#RkCCRL0CICMHRDO#CMCk8R##Cs3ERaH##RFOksCHRVDHCR#-
-RFbsPCH88MRFRRNMqQ1R1NRL#3H#RCaER Q  HR8#NODHRl#qRhYW)q)qYhaRu X)1 1R
m)-Q-RvQup Q7RhzBp7tQhRYqhR)Wq)aqhYwRmR)v Bh]qaQqApYQaR7qhRawQh1 1R)wmR z1
R--wRm)qqRu)BaQz)pqR)uzu m13ERaC#RkCFsRVER0CFR#kCsORDVHCER#NRDDHCM8lVMH$-
-R8NMRDEF8 RQ E RNDslCR##VlsFR$NMRl8NN#oCRRFsDLHNH0DH$sRNHM#HokRF0VRFRC0E
R--kR#C0sECC3FV

---a-RERH#b	NONRoClRN$LlCRFV8HHRC80HFRMkOD8NCR808HHNFMDNR80sNRCHJksRC8L0$RF#FD,-
-R0LkRRH0l0k#RRHMMIFRNO$REoNMCER0CGRC0MCsNHDRMs0CVCNO#sRFRl#Hk0DNHRFMLNCEPsHF
R--F0VRE8CRCs#OHHb0FRM3QH0R#CRbs#lH#DHLCFR0R8N8RlOFl0CM#MRN8s/FR0N0skHL0RC#0-F
-ER0CNRbOo	NCCR8OsDNNF0HMR#,LRk0MRF00OFREoNMCsRFRD8CCR0CNRM$FosHHDMNRMDHCF#RV-
-RC0ERObN	CNoRO8CDNNs0MHF3ERaCNRbOo	NCFRL8l$RNL$RCERONCMo8MRFDH$RMORNO8FsNCMO
R--IEH0RC0ERs0ClF#RV3R(4MRN83R(.VRFRH0E#0R#NNM8s
83---
-HRa0RDCRRRRR1:R08NMNRs8ep]7RM1$0#ECHu#RNNO	oRC#5 Q  0R18jR4(dn3-g4g(h,Rz)v QAB_Q
a2---
-HRpLssN$RRRRa:RERH#b	NONRoC#DENDCRLRlOFbCHD8MRH0NFRRLDHs$NsRl#$LHFDODND$-
-RRRRRRRRRRRR:NRMlRC8Q   3-
-
R--7CCPDCFbs:#RR Q  qR711BR$EM0C##HRsWF	oHMRFtsk
b3---
-kRus#bFCRRRRa:RERH#b	NONRoC8HCVMRC#MCklsRHO0C$b#MRN8sRNHl0ECO0HRMVkOF0HM-#
-RRRRRRRRRRRRV:RFksR#ICRHR0E#0$MEHC##FR0F3D#RFaIRlMkCOsHRb0$CN#Rs8CRCMVHC
8:-R-RRRRRRRRRRRR:->-RR1zhQ th7s:RCCbs#0CM#MRNR1zhQ th7kRMlsLCRRHMP0COFVsRF
sl-R-RRRRRRRRRRRR:->-RRt1Qh: 7RbsCsCC#MR0#NQR1t7h RlMkLRCsHPMRCFO0sFRVs-l
-RRRRRRRRRRRRa:RELCRNR#CClDCCRM00C$bRRH#0C$bRaAQ3-
-RRRRRRRRRRRR:ERaCCRDVF0l#L0RHH0R#sR0CCN08#RNRC0ER#lF0HR#oVMHHMON0HRL0-3
-RRRRRRRRRRRR1:RHCoM8CRPOs0F#sRNCCRsb#sCCCM08MRHRF0I'O#RFDlbCMlC0FRVs
l3-R-RRRRRRRRRRRR:a#EHRObN	CNoRMOF0MNH#PRFCFsDN88CRHNs0CEl0RHOFsbCNs0F#MRF
R--RRRRRRRRR:RRRC0ERt1QhR 7NRM8zQh1t7h Rb0$CR#3aRECb	NONRoCNFD#RMOF0MNH#-
-RRRRRRRRRRRR:#RkCDVkRb0$CFROMsPC#MHF#kRVMHO0F,M#RFODO8	RCO0C0MHF
R--RRRRRRRRR:RRRMVkOF0HMR#,NRM8FC0Es0RkH0DH$kRVMHO0F3M#
R--RRRRRRRRR:RR
R--RRRRRRRRR:RRRRQVNRM$Nksol0CMRR0FNkRVMHO0FHMR#RRNMDkDRsNsNR$,NkRMDNDRs$sNR
H#-R-RRRRRRRRRRRR:skC0s8MCRG5CO0CbH#FM,VRHR$NM,sRNCFRM0RC8HHM8PkH8N$DD2-3
--
-R0hFCRRRRRRR:FRhRO8CDNNs0MHF#sRFRV8CH0MHH#FMRN#EDLDRCMRHO8DkCH8RMF,Rs-
-RRRRRRRRRRRR:GRCO8DkCV8RsRFl0#EHRObN	CNo3ERaCbR"NNO	o8CRCNODsHN0FRM"8HCVM
C#-R-RRRRRRRRRRRR:0REC0C$b##,Rk$L0b,C#R8NMRO8CDNNs0MHF#VRFRvhz B)Q_aAQ3ERaC-
-RRRRRRRRRRRR:zRhvQ )BQ_AaNRbOo	NCFRL8#$REDNDRRLCO#FMHs8CC08REVCRFNslD-
-RRRRRRRRRRRR:CR8VHHM0MHFRRFV0REC#NClMO0H#VRFRH0E#NRbOo	NCa3RFRFD8CCPDCFbs-#
-RRRRRRRRRRRRl:RNO$RE#FFCFR0RbHlDCClM00REbCRNNO	oLCRFR8$H0MRElCRFR#0CHVVOMHC0-
-RRRRRRRRRRRR:NRlMsMCRNNPHLDND0CRFER0C
l3-R-RRRRRRRRRR
R:---R----------------------------------------------------------------------------
R--e#CsHRFMR:RRRc.3
R--7CN0RRRRR:RRRR4.qHbsDgR4g-6
--R--------------------------------------------------------------------------
--
ObN	CNoRvhz B)Q_aAQR
H#RFROMN#0MB0RF)b$H0oEhHF0ORC:1Qa)hRt
RRRRRR:="bBF$osHE�0RRg4g( RQ R 3qRDDsEHo0s#RCs#CP3C8"
;
R-R-============================================================================
-RR-kRhlHCsOsRqsRN$aC$bRV7CH0MHH#FM
-RR-============================================================================R

Rb0$ChRz1hQt H7R#sRNsRN$5ahqzp)qRMsNo<CR>RR2FAVRQ
a;R$R0b1CRQ th7#RHRsNsN5$Rhzqa)RqpsoNMC>R<RF2RVQRAa
;
R-R-============================================================================
-RR-sRqHl0ECO0HRCmbsFN0s
#:R-R-============================================================================
R
R-Q-R8q:R3R4
RMVkOF0HMNR"LR#"5tq):QR1t7h 2CRs0MksRt1Qh; 7RR--HLMRF
8$R-R-R#)CkRD0#0kL$:bCRt1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:)kC0sRM#0RECNFL#DCk0RDPNkFCRVRRN1hQt P7RCFO0s)Rqt
3
R-R-R:Q8R.q3
VRRk0MOHRFM"R-"5tq):QR1t7h 2CRs0MksRt1QhR 7=">RkH#lM"k#;R
R-)-RCD#k0kR#Lb0$C1:RQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CR)0Mks#ER0CNRPDRkCF0VREkCRM$NsRMlHkF#RbNCs0MHFRRFMNR
R-R-RRRRRR1RRQ th7CRPOs0FRtq)3R

R=--=========================================================================
==
-RR-8RQ:3RqdR
RVOkM0MHFR""+R,5pRR):zQh1t7h 2CRs0MksR1zhQ th7>R=RD"bk;#"
-RR-CR)#0kDRL#k0C$b:hRz1hQt v75qpX5'hp t,a]Rp)' aht]42-RI8FMR0FjR2
RR--)kC#DR0:q#88RF0IR1zhQ th7CRPOs0F#ER0Nl0RNL$RCVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RqcR
RVOkM0MHFR""+R,5pRR):1hQt R72skC0s1MRQ th7>R=Rb"#D"k#;R
R-)-RCD#k0kR#Lb0$C1:RQ th7q5vX'5ppt haR],) 'ph]ta2R-48MFI0jFR2R
R-)-RCD#k0q:R8R8#0RIF1hQt P7RCFO0s0#RERN0lRN$LFCRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8q:R3R6
RMVkOF0HM+R""pR5:hRz1hQt R7;)h:Rq)azqRp2skC0szMRht1QhR 7=">Rb#Dk"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0q:R8R8#NzMRht1QhR 7P0COFRs,pI,RHR0ENFRMMoMCNP0HChRQa  t)),R3R

RR--QR8:q
3nRkRVMHO0F"MR+5"Rph:Rq)azqRp;)z:Rht1Qh2 7R0sCkRsMzQh1t7h RR=>"kbD#
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:q#88RMNRFCMMoHN0PQCRhta  R),pI,RHR0ENzMRht1QhR 7P0COFRs,)
3
R-R-R:Q8R(q3
VRRk0MOHRFM"R+"5Rp:Q hat; )RR):1hQt R72skC0s1MRQ th7>R=Rb"#D"k#;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:q#88RRNMQ hat, )Rlp5NL$RCFRb#HH0PFCRsCRMoHN0P,C2RR0FNQR1t7h 
-RR-CRPOs0F,3R)
R
R-Q-R8q:R3RU
RMVkOF0HM+R""pR5:QR1t7h ;:R)RaQh )t 2CRs0MksRt1QhR 7=">R#kbD#
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:8Rq8N#RRt1QhR 7P0COFRs,p0,RFMRNRaQh )t ,3R)
R
R-=-==========================================================================
=
R-R-R:Q8Rgq3
VRRk0MOHRFM"R-"5Rp,)z:Rht1Qh2 7R0sCkRsMzQh1t7h RR=>"MlHk;#"
-RR-CR)#0kDRL#k0C$b:hRz1hQt v75qpX5'hp t,a]Rp)' aht]42-RI8FMR0FjR2
RR--)kC#DR0:10kLs0NO#IR0FhRz1hQt P7RCFO0s0#RERN0lRN$LFCRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8q:R3
4jRkRVMHO0F"MR-5"Rp),R:QR1t7h 2CRs0MksRt1QhR 7=">R#MlHk;#"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5Xvq5pp' aht]),R'hp t2a]-84RF0IMF2Rj
-RR-CR)#0kD:kR1LN0sOR0#NQR1t7h ROPC0,FsRR),VlsFRFNM0sECRt1QhR 7P0COFRs,pR,
RR--RRRRRRRR00ENR$lNR#bF#DHL$CRLRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R4q34R
RVOkM0MHFR""-R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMhRz1hQt =7R>lR"H#Mk"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k01:RksL0N#O0RMNRFCMMoHN0PQCRhta  R),)V,RsRFlNzMRht1QhR 7P0COFRs,p
3
R-R-R:Q8R4q3.R
RVOkM0MHFR""-R:5pRahqzp)q;:R)R1zhQ th7s2RCs0kMhRz1hQt =7R>lR"H#Mk"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RksL0N#O0RRNMzQh1t7h ROPC0,FsRR),VlsFRMNRFCMMoHN0PQCRhta  R),p
3
R-R-R:Q8R4q3dR
RVOkM0MHFR""-R:5pRt1Qh; 7RR):Q hat2 )R0sCkRsM1hQt =7R>#R"lkHM#
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:kR1LN0sOR0#NQMRhta  R),)V,RsRFlNQR1t7h ROPC0,FsR
p3
-RR-8RQ:3Rq4Rc
RMVkOF0HM-R""pR5:hRQa  t));R:QR1t7h 2CRs0MksRt1QhR 7=">R#MlHk;#"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RksL0N#O0R1NRQ th7CRPOs0F,,R)RFVslMRNRaQh )t ,3Rp
R
R-=-==========================================================================
=
R-R-R:Q8R4q36R
RVOkM0MHFR""*R,5pRR):zQh1t7h 2CRs0MksR1zhQ th7>R=Rk"lD;0"
-RR-CR)#0kDRL#k0C$b:hRz1hQt 575p 'ph]ta+p)' aht]2-4RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slRC0ERDlk0DHbH0ONHRFMFsbCNF0HMMRFRF0IR1zhQ th7CRPOs0F#R
R-R-RRRRRR0RRERN0lRN$b#F#H$LDRRLCF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:qn34
VRRk0MOHRFM"R*"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"k#lD;0"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5'5ppt ha)]+'hp t-a]482RF0IMF2Rj
-RR-CR)#0kD:kRvDb0HD#HCRF0IRt1QhR 7P0COFRs#00ENR$lNR#bF#DHL$CRLR
FVR-R-RRRRRRRRRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3Rq4R(
RMVkOF0HM*R""pR5:hRz1hQt R7;)h:Rq)azqRp2skC0szMRht1QhR 7=">Rl0kD"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5'5ppt hap]+'hp t-a]482RF0IMF2Rj
-RR-CR)#0kD:kRvDb0HD#HCRRNMzQh1t7h ROPC0,FsRRp,IEH0RMNRFCMMoHN0PRC
RR--RRRRRRRRQ hat, )RR)3)#RHRMOFP0CsC08RFMRNR1zhQ th7CRPOs0FR
FVR-R-RRRRRRRRRx#HC'Rppt haL]RCsVFCkRlDb0HDNHO0MHF3R

RR--QR8:qU34
VRRk0MOHRFM"R*"5Rp:hzqa);qpRR):zQh1t7h 2CRs0MksR1zhQ th7>R=Rk"lD;0"
-RR-CR)#0kDRL#k0C$b:hRz1hQt 575) 'ph]ta+p)' aht]2-4RI8FMR0FjR2
RR--)kC#DR0:v0kDHHbDCN#RMhRz1hQt P7RCFO0s),R,HRI0NERRMMFMNCo0CHP
-RR-RRRRRRRRhRQa  t)p,R3RRpHO#RFCMPs80CRR0FNzMRht1QhR 7P0COFFsRVR
R-R-RRRRRR#RRHRxC) 'ph]taRVLCFRsCl0kDHHbDOHN0F
M3
-RR-8RQ:3Rq4Rg
RMVkOF0HM*R""pR5:QR1t7h ;:R)RaQh )t 2CRs0MksRt1QhR 7=">R#Dlk0
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 75pp' aht]'+ppt ha4]-2FR8IFM0R
j2R-R-R#)Ck:D0RDvk0DHbHRC#NQR1t7h ROPC0,FsRRp,IEH0RRNMQ hat, )RR)3)#RH
-RR-RRRRRRRRFROMsPC0RC80NFRRt1QhR 7P0COFFsRVHR#xpCR'hp tRa]LFCVsRC
RR--RRRRRRRRl0kDHHbDOHN0F
M3
-RR-8RQ:3Rq.Rj
RMVkOF0HM*R""pR5:hRQa  t));R:QR1t7h 2CRs0MksRt1QhR 7=">R#Dlk0
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 75p)' aht]'+)pt ha4]-2FR8IFM0R
j2R-R-R#)Ck:D0RDvk0DHbHRC#NQR1t7h ROPC0,FsRR),IEH0RRNMQ hat, )RRp3p#RH
-RR-RRRRRRRRFROMsPC0RC80NFRRt1QhR 7P0COFFsRVHR#x)CR'hp tRa]LFCVsRC
RR--RRRRRRRRl0kDHHbDOHN0F
M3
-RR-============================================================================R
R-R-
RR--h ma:VRQRO#CFRM8Nksol0CMRRH#xFCsRsVFR""/RCFbsFN0sN,RRP#CC0sH$CRDP
CDR-R-RRRRRFRRV)R )Rm)HH#R#C#k8
3
R-R-R:Q8R.q34R
RVOkM0MHFR""/R,5pRR):zQh1t7h 2CRs0MksR1zhQ th7>R=RH"8P
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#NzMRht1QhR 7P0COFRs,pL,R$MRNFC0EshRz1hQt P7RCFO0s),R3R

RR--QR8:q.3.
VRRk0MOHRFM"R/"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"P8H"R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RP7HH#8CRRNM1hQt P7RCFO0sp,R,$RLRFNM0sECRt1QhR 7P0COFRs,)
3
R-R-R:Q8R.q3dR
RVOkM0MHFR""/R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMhRz1hQt =7R>8R"H;P"
-RR-CR)#0kDRL#k0C$b:hRz1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RP7HH#8CRRNMzQh1t7h ROPC0,FsRRp,LN$RRMMFMNCo0CHPRaQh )t ,3R)
-RR-RRRRRRRRVRQR_hmmAw_Q5a1)>2RRpp' aht]s,RCD#k0#RHRk0sM0ONC08RF'Rppt ha
]3
-RR-8RQ:3Rq.Rc
RMVkOF0HM/R""pR5:qRhaqz)p);R:hRz1hQt R72skC0szMRht1QhR 7=">RMH#8P
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#NFRMMoMCNP0HChRQa  t)p,R,$RLRRNMzQh1t7h ROPC0,FsR
)3R-R-RRRRRRRRRRQVhmm_wQ_Aap152RR>) 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rp)' aht]
3
R-R-R:Q8R.q36R
RVOkM0MHFR""/R:5pRt1Qh; 7RR):Q hat2 )R0sCkRsM1hQt =7R>MR"#H#8P
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#RRN1hQt P7RCFO0sp,R,$RLRRNMQ hat, )R
)3R-R-RRRRRRRRRRQVhmm_wQ_Aa)152RR>p 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rpp' aht]
3
R-R-R:Q8R.q3nR
RVOkM0MHFR""/R:5pRaQh )t ;:R)Rt1Qh2 7R0sCkRsM1hQt =7R>MR"#H#8P
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#MRNRaQh )t ,,RpRRL$NQR1t7h ROPC0,FsR
)3R-R-RRRRRRRRRRQVhmm_wQ_Aap152RR>) 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rp)' aht]
3
R-R-============================================================================
-RR-R
R-h-Rm:a RRQV#FCOMN8RslokCRM0Hx#RCRsFVRFs"lsC"bRFC0sNFRs,NCR#PHCs0D$RCDPC
-RR-RRRRRRRF VR)))mRRH#Hk##C
83
-RR-8RQ:3Rq.R(
RMVkOF0HMsR"CRl"5Rp,)z:Rht1Qh2 7R0sCkRsMzQh1t7h RR=>"sM#C;l"
-RR-CR)#0kDRL#k0C$b:hRz1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"RlsCRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0s
#3
-RR-8RQ:3Rq.RU
RMVkOF0HMsR"CRl"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"#M#s"Cl;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRNpRM)8RRCNsRt1QhR 7P0COF3s#
R
R-Q-R8q:R3
.gRkRVMHO0F"MRs"ClR:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMhRz1hQt =7R>sR"C;l"
-RR-CR)#0kDRL#k0C$b:hRz1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"RlsCRR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8RR)HN#R
-RR-RRRRRRRRFRMMoMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:qj3d
VRRk0MOHRFM"lsC"pR5:qRhaqz)p);R:hRz1hQt R72skC0szMRht1QhR 7=">RMC#sl
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRH)R#MRNR1zhQ th7CRPOs0FR8NMRHpR#
RNR-R-RRRRRRRRRMMFMNCo0CHPRaQh )t 3R
R-Q-RVmRh__mwA1Qa5Rp2>'R)pt haR],skC#DH0R#sR0kNMO0RC80)FR'hp t3a]
R
R-Q-R8q:R3
d4RkRVMHO0F"MRs"ClR:5pRt1Qh; 7RR):Q hat2 )R0sCkRsM1hQt =7R>MR"#C#sl
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpCRsl"R)RCIEspCRRRH#1hQt P7RCFO0sMRN8RR)HN#RMhRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:q.3d
VRRk0MOHRFM"lsC"pR5:hRQa  t));R:QR1t7h 2CRs0MksRt1QhR 7=">RMs##C;l"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsC)#RHRt1QhR 7P0COFNsRMp8RRRH#NQMRhta  
)3R-R-RRRRRRRRRRQVhmm_wQ_Aap152RR>) 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rp)' aht]
3

-RR-============================================================================R
R-R-
RR--h ma:VRQRO#CFRM8Nksol0CMRRH#xFCsRsVFRF"l8F"RbNCs0,FsR#NRCsPCHR0$DCCPDR
R-R-RRRRRRRFV m)))#RHR#H#k3C8
R
R-Q-R8q:R3
ddRkRVMHO0F"MRl"F8R,5pRR):zQh1t7h 2CRs0MksR1zhQ th7>R=R#"Ml"F8;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpFRl8"R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COF3s#
R
R-Q-R8q:R3
dcRkRVMHO0F"MRl"F8R,5pRR):1hQt R72skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"R8lFRR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#Fs3R

RR--QR8:q63d
VRRk0MOHRFM"8lF"pR5:hRz1hQt R7;)h:Rq)azqRp2skC0szMRht1QhR 7=">Rl"F8;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpFRl8"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRM)8R
-RR-RRRRRRRR#RHRMNRFCMMoHN0PQCRhta  
)3R-R-RRRRRRRRRRQVhmm_wQ_Aa)152RR>p 'ph]ta,CRs#0kDRRH#0MskOCN08FR0Rpp' aht]
3
R-R-R:Q8Rdq3nR
RVOkM0MHFRF"l85"Rph:Rq)azqRp;)z:Rht1Qh2 7R0sCkRsMzQh1t7h RR=>"lM#F;8"
-RR-CR)#0kDRL#k0C$b:hRz1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"R8lFRR)"IsECCRR)HN#RMhRz1hQt P7RCFO0sMRN8
RpR-R-RRRRRRRRRRH#NFRMMoMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]R#sCkRD0H0#RsOkMN80CRR0F) 'ph]ta3R

RR--QR8:q(3d
VRRk0MOHRFM"8lF"pR5:QR1t7h ;:R)RaQh )t 2CRs0MksRt1QhR 7=">RMF#l8
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpFRl8"R)RCIEspCRRRH#NQR1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R
R-R-RRRRRRQRRVmRh__mwA1Qa5R)2>'Rppt haR],skC#DH0R#sR0kNMO0RC80pFR'hp t3a]
R
R-Q-R8q:R3
dURkRVMHO0F"MRl"F8R:5pRaQh )t ;:R)Rt1Qh2 7R0sCkRsM1hQt =7R>MR"#8lF"R;
RR--)kC#D#0Rk$L0bRC:1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RlBFbCk0#pR"R8lFRR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NQR1t7h ROPC03Fs
-RR-RRRRRRRRVRQR_hmmAw_Q5a1p>2RRp)' aht]s,RCD#k0#RHRk0sM0ONC08RF'R)pt ha
]3
-
-============================================================================
-RR-8RQ:3RqdRg
RMVkOF0HMHRVMD8_ClV0FR#05tq)Rz:Rht1Qh; 7R:YRRaAQ2CRs0MksRaQh )t ;R
R-)-RCD#k0kR#Lb0$CQ:Rhta  R)
RR--)kC#DR0:w8HM#ER0CCRDVF0l#F0ROsOksOCMCVRFRC0ERDPNkFCRVRRYHqMR)
t3R-R-RRRRRRRRR0)Ck#sMRC0ER8HMCFGRVER0CORFOsksCCMORRHVHC0RG0H##F,Rs4R-REF0CHsI#
C3
-RR-8RQ:3RqcRj
RMVkOF0HMHRVMD8_ClV0FR#05tq)R1:RQ th7Y;RRA:RQRa2skC0sQMRhta  
);R-R-R#)CkRD0#0kL$:bCRaQh )t 
-RR-CR)#0kD:HRwMR8#0RECD0CVl0F#ROFOkCssMROCF0VREPCRNCDkRRFVYMRHRtq)3R
R-R-RRRRRR)RRCs0kM0#REHCRMG8CRRFV0RECFkOOsMsCOHCRV0RHRHCG#,0#RRFs-F4R0sECICH#3R

RR--QR8:q43c
VRRk0MOHRFMV8HM_osHEF0l#50RqR)t:hRz1hQt R7;YRR:A2QaR0sCkRsMQ hat; )
-RR-CR)#0kDRL#k0C$b:hRQa  t)R
R-)-RCD#k0w:RH#M8RC0ERVDC0#lF0ORFOsksCCMORRFV0RECPkNDCVRFRHYRM)RqtR3
RR--RRRRRRRR)kC0sRM#0RECHCM8GVRFRC0EROFOkCssMROCHHVR0GRCH##0,sRFRR-4FC0Es#IHC
3
R-R-R:Q8Rcq3.R
RVOkM0MHFRMVH8H_solE0FR#05tq)R1:RQ th7Y;RRA:RQRa2skC0sQMRhta  
);R-R-R#)CkRD0#0kL$:bCRaQh )t 
-RR-CR)#0kD:HRwMR8#0RECD0CVl0F#ROFOkCssMROCF0VREPCRNCDkRRFVYMRHRtq)3R
R-R-RRRRRR)RRCs0kM0#REHCRMG8CRRFV0RECFkOOsMsCOHCRV0RHRHCG#,0#RRFs-F4R0sECICH#3


R-R-============================================================================
-RR-FRBlsbNHM#FRCmbsFN0sR#
R=--=========================================================================
==
-RR-8RQ:3RB4R
RVOkM0MHFR"">R,5pRR):zQh1t7h 2CRs0MksRmAmph qRR=>"0ko"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3R.
RMVkOF0HM>R""pR5,:R)Rt1Qh2 7R0sCkRsMApmm Rqh=">R#"o0;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRR8NMRN)Rs1CRQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B
3dRkRVMHO0F"MR>5"Rph:Rq)azqRp;)z:Rht1Qh2 7R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRMMFMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8RcB3
VRRk0MOHRFM"R>"5Rp:Q hat; )RR):1hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#RRNQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R6B3
VRRk0MOHRFM"R>"5Rp:zQh1t7h ;:R)Rahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-8RQ:3RBnR
RVOkM0MHFR"">R:5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRQNRhta  
)3
-RR-============================================================================R

RR--QR8:B
3(RkRVMHO0F"MR<5"Rp),R:hRz1hQt R72skC0sAMRm mpq=hR>kR"D;0"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RUB3
VRRk0MOHRFM"R<"5Rp,)1:RQ th7s2RCs0kMmRAmqp h>R=RD"#0
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRNpRM)8RRCNsRt1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBgR
RVOkM0MHFR""<R:5pRahqzp)q;:R)R1zhQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRMNRFCMMoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
4jRkRVMHO0F"MR<5"RpQ:Rhta  R);)1:RQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R4B34R
RVOkM0MHFR""<R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
4.RkRVMHO0F"MR<5"Rp1:RQ th7);R:hRQa  t)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHR1NRQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RMhRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3
4dRkRVMHO0F"MR<R="5Rp,)z:Rht1Qh2 7R0sCkRsMApmm Rqh=">Rk"DC;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
4cRkRVMHO0F"MR<R="5Rp,)1:RQ th7s2RCs0kMmRAmqp h>R=RD"#C
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
46RkRVMHO0F"MR<R="5Rp:hzqa);qpRR):zQh1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRMNRFCMMoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
4nRkRVMHO0F"MR<R="5Rp:Q hat; )RR):1hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NQR1t7h ROPC03Fs
R
R-Q-R8B:R3
4(RkRVMHO0F"MR<R="5Rp:zQh1t7h ;:R)Rahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
4URkRVMHO0F"MR<R="5Rp:1hQt R7;)Q:Rhta  R)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R4B3gR
RVOkM0MHFR=">"pR5,:R)R1zhQ th7s2RCs0kMmRAmqp h>R=Ro"kC
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R.B3jR
RVOkM0MHFR=">"pR5,:R)Rt1Qh2 7R0sCkRsMApmm Rqh=">R#"oC;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R.B34R
RVOkM0MHFR=">"pR5:qRhaqz)p);R:hRz1hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRMMFMNCo0CHPRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz1hQt P7RCFO0s
3
R-R-R:Q8R.B3.R
RVOkM0MHFR=">"pR5:hRQa  t));R:QR1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R.B3dR
RVOkM0MHFR=">"pR5:hRz1hQt R7;)h:Rq)azqRp2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMoMCNP0HChRQa  t)
3
R-R-R:Q8R.B3cR
RVOkM0MHFR=">"pR5:QR1t7h ;:R)RaQh )t 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCp#RHR1NRQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RMhRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3
.6RkRVMHO0F"MR=5"Rp),R:hRz1hQt R72skC0sAMRm mpq=hR>CR"J
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bn3.
VRRk0MOHRFM"R="5Rp,)1:RQ th7s2RCs0kMmRAmqp h>R=RJ"C"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R.B3(R
RVOkM0MHFR""=R:5pRahqzp)q;:R)R1zhQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRMNRFCMMoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
.URkRVMHO0F"MR=5"RpQ:Rhta  R);)1:RQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R.B3gR
RVOkM0MHFR""=R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
djRkRVMHO0F"MR=5"Rp1:RQ th7);R:hRQa  t)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHR1NRQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RMhRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3
d4RkRVMHO0F"MR/R="5Rp,)z:Rht1Qh2 7R0sCkRsMApmm Rqh=">RMCF0J
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RdB3.R
RVOkM0MHFR="/"pR5,:R)Rt1Qh2 7R0sCkRsMApmm Rqh=">RMCF0J
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
ddRkRVMHO0F"MR/R="5Rp:hzqa);qpRR):zQh1t7h 2CRs0MksRmAmph qRR=>"0MFC;J"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBdRc
RMVkOF0HM/R"=5"RpQ:Rhta  R);)1:RQ th7s2RCs0kMmRAmqp h>R=RF"M0"CJ;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8RdB36R
RVOkM0MHFR="/"pR5:hRz1hQt R7;)h:Rq)azqRp2skC0sAMRm mpq=hR>MR"FJ0C"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

RR--QR8:Bn3d
VRRk0MOHRFM""/=R:5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm Rqh=">RMCF0J
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
-
-R:Q8RdB3(R
RVOkM0MHFRhvQQvvzR,5pR:)RR1zhQ th7s2RCs0kMhRz1hQt 
7;R-R-R#)CkRD0#0kL$:bCR1zhQ th7R
R-)-RCD#k0):RCs0kM0#REDCRCC##sVRFRF0IR1zhQ th7CRPOs0F#ER0Nl0RNL$RCR
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
dURkRVMHO0FvMRQvhQz5vRp),RR1:RQ th7s2RCs0kMQR1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7R
R-)-RCD#k0):RCs0kM0#REDCRCC##sVRFRF0IRt1QhR 7P0COFRs#00ENR$lNR
LCR-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RdB3gR
RVOkM0MHFRhvQQvvzRR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRRMMFMNCo0CHPRaQh )t ,,RpR8NM
-RR-RRRRRRRRMRNR1zhQ th7CRPOs0F,3R)
R
R-Q-R8B:R3
cjRkRVMHO0FvMRQvhQz5vRpRR:Q hat; )R:)RRt1Qh2 7R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRMhRQa  t)p,R,MRN8RRN1hQt R7
RR--RRRRRRRRP0COFRs,)
3
R-R-R:Q8RcB34R
RVOkM0MHFRhvQQvvzRR5p:hRz1hQt R7;)RR:hzqa)2qpR0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRMhRz1hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRRMMFMNCo0CHPRaQh )t ,3R)
R
R-Q-R8B:R3
c.RkRVMHO0FvMRQvhQz5vRpRR:1hQt R7;)RR:Q hat2 )R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRRt1QhR 7P0COFRs,pN,RMR8
RR--RRRRRRRRNQMRhta  R),)
3
R-R-============================================================================
R
R-Q-R8B:R3
cdRkRVMHO0FvMRqvXQz5vRp),RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ERCosNs0CRRFV0RIFzQh1t7h ROPC0#FsRN0E0NRl$CRL
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBcRc
RMVkOF0HMqRvXzQvvpR5,RR):QR1t7h 2CRs0MksRt1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 
-RR-CR)#0kD:CR)0Mks#ER0CsRoCCN0sVRFRF0IRt1QhR 7P0COFRs#00ENR$lNR
LCR-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RcB36R
RVOkM0MHFRXvqQvvzRR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ERCosNs0CRRFVNFRMMoMCNP0HChRQa  t)p,R,MRN8R
R-R-RRRRRRNRRMhRz1hQt P7RCFO0s),R3R

RR--QR8:Bn3c
VRRk0MOHRFMvQqXvRzv5:pRRaQh )t ;RR):QR1t7h 2CRs0MksRt1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 
-RR-CR)#0kD:CR)0Mks#ER0CsRoCCN0sVRFRRNMQ hat, )RRp,NRM8NQR1t7h 
-RR-RRRRRRRRCRPOs0F,3R)
R
R-Q-R8B:R3
c(RkRVMHO0FvMRqvXQz5vRpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMhRz1hQt 
7;R-R-R#)CkRD0#0kL$:bCR1zhQ th7R
R-)-RCD#k0):RCs0kM0#REoCRs0CNCFsRVMRNR1zhQ th7CRPOs0F,,RpR8NM
-RR-RRRRRRRRRRNMMFMC0oNHRPCQ hat, )R
)3
-RR-8RQ:3RBcRU
RMVkOF0HMqRvXzQvvpR5R1:RQ th7);RRQ:Rhta  R)2skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt R7
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsFNVRRt1QhR 7P0COFRs,pN,RMR8
RR--RRRRRRRRNQMRhta  R),)
3
R-R-============================================================================
R
R-Q-R8B:R3
cgRkRVMHO0F"MR?R>"5Rp,)RR:zQh1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB6Rj
RMVkOF0HM?R">5"Rp),RR1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R6B34R
RVOkM0MHFR>"?"pR5Rh:Rq)azqRp;)RR:zQh1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB6R.
RMVkOF0HM?R">5"RpRR:Q hat; )R:)RRt1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RRt1QhR 7P0COF
s3
-RR-8RQ:3RB6Rd
RMVkOF0HM?R">5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
6cRkRVMHO0F"MR?R>"5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NQR1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R6B36R
RVOkM0MHFR<"?"pR5,RR):hRz1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bn36
VRRk0MOHRFM""?<R,5pR:)RRt1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
6(RkRVMHO0F"MR?R<"5:pRRahqzp)q;RR):hRz1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:BU36
VRRk0MOHRFM""?<RR5p:hRQa  t));RR1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R6B3gR
RVOkM0MHFR<"?"pR5Rz:Rht1Qh; 7R:)RRahqzp)q2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-8RQ:3RBnRj
RMVkOF0HM?R"<5"RpRR:1hQt R7;)RR:Q hat2 )R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8RnB34R
RVOkM0MHFR<"?=5"Rp),RRz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBnR.
RMVkOF0HM?R"<R="5Rp,)RR:1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
ndRkRVMHO0F"MR?"<=RR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBnRc
RMVkOF0HM?R"<R="5:pRRaQh )t ;RR):QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8RnB36R
RVOkM0MHFR<"?=5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

RR--QR8:Bn3n
VRRk0MOHRFM"=?<"pR5R1:RQ th7);RRQ:Rhta  R)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8RnB3(R
RVOkM0MHFR>"?=5"Rp),RRz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBnRU
RMVkOF0HM?R">R="5Rp,)RR:1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
ngRkRVMHO0F"MR?">=RR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB(Rj
RMVkOF0HM?R">R="5:pRRaQh )t ;RR):QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R(B34R
RVOkM0MHFR>"?=5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

RR--QR8:B.3(
VRRk0MOHRFM"=?>"pR5R1:RQ th7);RRQ:Rhta  R)2skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
R
R-=-==========================================================================
=
R-R-R:Q8R(B3dR
RVOkM0MHFR="?"pR5,RR):hRz1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bc3(
VRRk0MOHRFM""?=R,5pR:)RRt1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAaR
R-)-RCD#k0B:RFklb0RC#"=pRRR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
(6RkRVMHO0F"MR?R="5:pRRahqzp)q;RR):hRz1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:Bn3(
VRRk0MOHRFM""?=RR5p:hRQa  t));RR1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNRt1QhR 7P0COF
s3
-RR-8RQ:3RB(R(
RMVkOF0HM?R"=5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
(URkRVMHO0F"MR?R="5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#N1MRQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RMhRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3
(gRkRVMHO0F"MR?"/=R,5pR:)RR1zhQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRNpRM)8RRCNsR1zhQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bj3U
VRRk0MOHRFM"=?/"pR5,RR):QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RUB34R
RVOkM0MHFR/"?=5"RpRR:hzqa);qpR:)RR1zhQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:B.3U
VRRk0MOHRFM"=?/"pR5RQ:Rhta  R);)RR:1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#N1MRQ th7CRPOs0F3R

RR--QR8:Bd3U
VRRk0MOHRFM"=?/"pR5Rz:Rht1Qh; 7R:)RRahqzp)q2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
UcRkRVMHO0F"MR?"/=RR5p:QR1t7h ;RR):hRQa  t)s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A
QaR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#MRNRt1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRRNMQ hat3 )
R

R=--=========================================================================
==R-R-RH1EVN0RM)8RF00NCkRwMHO0F
M#R-R-============================================================================
R
R-Q-R81:R3R4
RMVkOF0HM]R1Q_wapa wR)5qtz:Rht1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsMzQh1t7h RR=>"D#D"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRN#VEH0C-DVF0RMMRNR1zhQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0R0AHR''j3R
R-R-RRRRRRaRREBCRmazhRVDC0#lF0HRL0N#RsDCRF3#0
R
R-Q-R81:R3R.
RMVkOF0HM]R1Q_wa)]QtaqR5)Rt:zQh1t7h ;mRBz:haRahqzp)q2CRs0MksR1zhQ th7>R=Rs"#D
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRussVFlN#RRH#EVs0-H0oERRFMNzMRht1QhR 7P0COFBsRmazhRl0HC
#3R-R-RRRRRRRRRCaEROPNN80CR#bFHF0HMN#RsVCRHCDD8HRI0AERH'0Rj
'3R-R-RRRRRRRRRCaERzBmhsaRH0oEl0F#R0LH#sRNCFRD#
03
-RR-8RQ:3R1dR
RVOkM0MHFRQ1]wpa_ Rwa5tq):QR1t7h ;mRBz:haRahqzp)q2CRs0MksRt1QhR 7=">R#"DD;R
R-)-RCD#k0kR#Lb0$C1:RQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRussVFlN#RRH#EVD0-CRV0FNMRRt1QhR 7P0COFBsRmazhRl0HC
#3R-R-RRRRRRRRRCaEROPNN80CR#bFHF0HMN#RsVCRHCDD8HRI0AERH'0Rj
'3R-R-RRRRRRRRRCaERzBmhDaRClV0FR#0L#H0RCNsR#DF0
3
R-R-R:Q8Rc13
VRRk0MOHRFM1w]QaQ_)tR]a5tq):QR1t7h ;mRBz:haRahqzp)q2CRs0MksRt1QhR 7=">R#"sN;R
R-)-RCD#k0kR#Lb0$C1:RQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRussVFlN#RRH#EVs0-H0oERRFMNQR1t7h ROPC0RFsBhmzaHR0l3C#
-RR-RRRRRRRRERaCNRPOCN08FRb#HH0FRM#NRsCVDHDCI8RHR0E0RECD0CVl0F#R0LH,)Rqt 'pw
a3R-R-RRRRRRRRRCaERzBmhsaRH0oEl0F#R0LH#sRNCFRD#
03
-RR-============================================================================R

RR--QR8:1
36RkRVMHO0F)MRmaaq  _pw5aRq:)tR1zhQ th7B;Rmazh:qRhaqz)ps2RCs0kMhRz1hQt =7R>sR"F;D"
-RR-CR)#0kDRL#k0C$b:hRz1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NFRs0CN0-VDC0VRFRRNMzQh1t7h ROPC0RFsBhmzaHR0l3C#
R
R-Q-R81:R3Rn
RMVkOF0HMmR)a qa_t)Q]5aRq:)tR1zhQ th7B;Rmazh:qRhaqz)ps2RCs0kMhRz1hQt =7R>sR"F;s"
-RR-CR)#0kDRL#k0C$b:hRz1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NFRs0CN0-osHEF0RVMRNR1zhQ th7CRPOs0FRzBmh0aRH#lC3R

RR--QR8:1
3(RkRVMHO0F)MRmaaq  _pw5aRq:)tRt1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsM1hQt =7R>sR"F;D"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRNDHFoORNDsNF00DC-CRV0FNVRRt1QhR 7P0COFBsRmazhRl0HC
#3
-RR-8RQ:3R1UR
RVOkM0MHFRa)mq_a )]QtaqR5)Rt:1hQt R7;Bhmzah:Rq)azqRp2skC0s1MRQ th7>R=RF"ss
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slRDNRFOoHNsDRF00NCH-soRE0FNVRRt1QhR 7P0COFBsRmazhRl0HC
#3
-RR-============================================================================R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1R3gHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1
3gRkRVMHO0F"MR#"DDR)5qtz:Rht1Qh; 7RzBmhRa:Q hat2 )R0sCkRsMzQh1t7h RR=>"D#D"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]wpa_ 5waq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14HjR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4jRkRVMHO0F"MR#"DDR)5qt1:RQ th7B;Rmazh:hRQa  t)s2RCs0kMQR1t7h RR=>"D#D"R;
RR--)kC#D#0Rk$L0bRC:1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_wp a)5qtB,Rmazh2R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1434RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R4134R
RVOkM0MHFRs"#D5"Rq:)tR1zhQ th7B;Rmazh:hRQa  t)s2RCs0kMhRz1hQt =7R>#R"s;D"
-RR-CR)#0kDRL#k0C$b:hRz1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_t)Q]qa5)Rt,Bhmza
2
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413.#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14R.
RMVkOF0HM#R"sRD"5tq):QR1t7h ;mRBz:haRaQh )t 2CRs0MksRt1QhR 7=">R#"sD;R
R-)-RCD#k0kR#Lb0$C1:RQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:QR1t7h 5Q1]w)a_Qat]51zhQ th7)5qtR2,Bhmza
22
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14HdR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4dRkRVMHO0F"MRs"FDR)5qtz:Rht1Qh; 7RzBmhRa:Q hat2 )R0sCkRsMzQh1t7h RR=>"DsF"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a pa w5tq),mRBz2ha
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0F1MR3R4cHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1c34
VRRk0MOHRFM"DsF"qR5)Rt:1hQt R7;BhmzaQ:Rhta  R)2skC0s1MRQ th7>R=RF"sD
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:)qmaap _ 5waq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14H6R#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
46RkRVMHO0F"MRs"FsR)5qtz:Rht1Qh; 7RzBmhRa:Q hat2 )R0sCkRsMzQh1t7h RR=>"ssF"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a )]Qta)5qtB,Rmazh2R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1n34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413nR
RVOkM0MHFRF"ss5"Rq:)tRt1Qh; 7RzBmhRa:Q hat2 )R0sCkRsM1hQt =7R>sR"F;s"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a )]Qta)5qtB,Rmazh2R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1(34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413(R
RVOkM0MHFRD"#N5"RqR)t:hRz1hQt R7;BhmzaRR:Q hat2 )R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]Qa _pwqa5)Rt,Bhmza
2
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413U#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14RU
RMVkOF0HM#R"DRN"5tq)R1:RQ th7B;RmazhRQ:Rhta  R)2skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_wp a)5qtB,Rmazh2R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1g34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413gR
RVOkM0MHFRs"#N5"RqR)t:hRz1hQt R7;BhmzaRR:Q hat2 )R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]QaQ_)t5]aq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R1.HjR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
.jRkRVMHO0F"MR#"sNR)5qtRR:1hQt R7;BhmzaRR:Q hat2 )R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]QaQ_)t5]aq,)tRzBmh
a2
R
R-=-==========================================================================R=
RR--)Q 1Zw Rk0MOH#FM
-RR-============================================================================R

RR--QR8:)
34RkRVMHO0F)MR Z1Q qR5)Rt:1hQt R7;h_ W1 QZ:qRhaqz)ps2RCs0kMQR1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7 5hWQ_1Z4 -RI8FMR0FjR2
RR--)kC#DR0:)HC#xRC#0REC1hQt P7RCFO0s)RqtFR0RC0ERC#bOHHVC#8RH3xC
-RR-RRRRRRRRFRaRCOsNR0CNNRDssoCROPC0,FsRC0ERIMCRCrDVF0l#R09LRH0bHF#0MHF#R
R-R-RRRRRRNRRsVCRHCDD8HRI00ERE#CRHRoMLRH05tq)'wp aR23WMECRk0sM0ONH,Mo
-RR-RRRRRRRRER0CHR#oLMRHH0R#CRs0MNHCN8RDoFMR0IHEER0CHRsolE0FR#0b0Ns3R

RR--QR8:)
3.RkRVMHO0F)MR Z1Q qR5)Rt:zQh1t7h ; RhWQ_1ZR :hzqa)2qpR0sCkRsMzQh1t7h RR=>"H0sl
";R-R-R#)CkRD0#0kL$:bCR1zhQ th7 5hWQ_1Z4 -RI8FMR0FjR2
RR--)kC#DR0:)HC#xRC#0RECzQh1t7h ROPC0RFsqR)t00FRE#CRbHCOV8HCRx#HCR3
RR--RRRRRRRRaOFRs0CNCRRNDoNsCPsRCFO0s0,REMCRCrIRD0CVl0F#9HRL0FRb#HH0F
M#R-R-RRRRRRRRRCNsRDVHDRC8IEH0R''j3ERWC0MRsOkMNM0Ho0,REDCRClV0FR#0L#H0
-RR-RRRRRRRRsRNCsR8FCbb8
3
RkRVMHO0F)MR Z1Q qR5)Rt,1 QZ_1) Rz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt 57R1 QZ_1) 'MDCo-0E4FR8IFM0R
j2
VRRk0MOHRFM)Q 1Z5 Rq,)tRZ1Q  _)1RR:1hQt R72skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th71R5Q_Z )' 1DoCM04E-RI8FMR0Fj
2

-RR-============================================================================R
R-B-RFCMPsF#HMkRwMHO0F
M#R-R-============================================================================
R
R-Q-R87:R3R4
RMVkOF0HMmRa_aQh )t R)5qtz:Rht1Qh2 7R0sCkRsMhzqa)Rqp=">RLHkV"R;
RR--)kC#D#0Rk$L0bRC:hzqa)3qpRDeNkOCRNFMM0CRLRoMCNP0HCHR#MROCbNNslCC0s#RHR
NMR-R-RRRRRRRRR1zhQ th7CRPOs0F3R
R-)-RCD#k0B:RFCMPsR0#0RECzQh1t7h ROPC0RFs0NFRMhRQa  t)
3
R-R-R:Q8R.73
VRRk0MOHRFMaQm_hta  5)Rq:)tRt1Qh2 7R0sCkRsMQ hatR )=">RL#kVH
";R-R-R#)CkRD0#0kL$:bCRaQh )t 
-RR-CR)#0kD:FRBMsPC0N#RRt1QhR 7P0COF0sRFMRNRaQh )t 3R

RR--QR8:7
3dRkRVMHO0FaMRmh_z1hQt 57Rq,)tRZ1Q h:Rq)azqRp2skC0szMRht1QhR 7=">R0lsH"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5Z1Q R-48MFI0jFR2R
R-)-RCD#k0B:RFCMPsR0#NFRMMoMCNP0HChRQa  t)FR0RRNMzQh1t7h ROPC0RFsIEH0
-RR-RRRRRRRRER0CbR#CVOHHRC8#CHx3R

RR--QR8:7
3cRkRVMHO0FaMRmQ_1t7h R)5qtQ:Rhta  R);1 QZ:qRhaqz)ps2RCs0kMQR1t7h RR=>"s#0H;l"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5Z1Q R-48MFI0jFR2R
R-)-RCD#k0B:RFCMPsR0#NQMRhta  0)RFRRN1hQt P7RCFO0sVRFRC0ERC#bOHHVC#8RH3xC
R
RVOkM0MHFR_amzQh1t7h R)5qtRR:hzqa);qpRZ1Q  _)1RR:zQh1t7h 2CRs0MksR1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 71 QZ_1) 'MDCo-0E4FR8IFM0R
j2
VRRk0MOHRFMa1m_Q th7qR5):tRRaQh )t ;QR1Z) _ :1RRt1Qh2 7R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt 175Q_Z )' 1DoCM04E-RI8FMR0Fj
2

-RR-============================================================================R
R-p-RFOoHNmDRbNCs0#Fs
-RR-============================================================================R

RR--QR8:p
34RkRVMHO0F"MRM"F0R:5pR1zhQ th7s2RCs0kMhRz1hQt =7R>MR"F;0"
-RR-CR)#0kDRL#k0C$b:hRz1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsaCl#IHCMRHP#CsH
FM
-RR-8RQ:3Rp.R
RVOkM0MHFRM"N85"Rp),R:hRz1hQt R72skC0szMRht1QhR 7=">RN"M8;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0FR7qhRCFbsHN0F
M
R-R-R:Q8Rdp3
VRRk0MOHRFM""FsR,5pRR):zQh1t7h 2CRs0MksR1zhQ th7>R=Rs"F"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0s)RmRCFbsHN0F
M
R-R-R:Q8Rcp3
VRRk0MOHRFM"MMN85"Rp),R:hRz1hQt R72skC0szMRht1QhR 7=">RM8NM"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sqRhhF7RbNCs0MHF
R
R-Q-R8p:R3R6
RMVkOF0HMMR"FRs"5Rp,)z:Rht1Qh2 7R0sCkRsMzQh1t7h RR=>"sMF"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0smRh)bRFC0sNH
FM
-RR-8RQ:3RpnR
RVOkM0MHFRF"Gs5"Rp),R:hRz1hQt R72skC0szMRht1QhR 7=">RG"Fs;R
R-)-RCD#k0kR#Lb0$Cz:Rht1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0FR)XmRCFbsHN0F
M
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR(p3RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R(p3
VRRk0MOHRFM"FGMs5"Rp),R:hRz1hQt R72skC0szMRht1QhR 7=">RGsMF"R;
RR--)kC#D#0Rk$L0bRC:zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0shRXmF)RbNCs0MHF
R
R-Q-R8p:R3RU
RMVkOF0HMMR"FR0"5Rp:1hQt R72skC0s1MRQ th7>R=RF"M0
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CRasHlI#HCRMsPC#MHF
R
R-Q-R8p:R3Rg
RMVkOF0HMNR"MR8"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"8NM"R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0RFsqRh7FsbCNF0HMR

RR--QR8:pj34
VRRk0MOHRFM""FsR,5pRR):1hQt R72skC0s1MRQ th7>R=Rs"F"R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0RFsmF)RbNCs0MHF
R
R-Q-R8p:R3
44RkRVMHO0F"MRM8NM"pR5,:R)Rt1Qh2 7R0sCkRsM1hQt =7R>MR"N"M8;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COFhsRqRh7FsbCNF0HMR

RR--QR8:p.34
VRRk0MOHRFM"sMF"pR5,:R)Rt1Qh2 7R0sCkRsM1hQt =7R>MR"F;s"
-RR-CR)#0kDRL#k0C$b:QR1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0smRh)bRFC0sNH
FM
-RR-8RQ:3Rp4Rd
RMVkOF0HMGR"FRs"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"sGF"R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0RFsXRm)FsbCNF0HMR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpc34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R4p3cR
RVOkM0MHFRM"GFRs"5Rp,)1:RQ th7s2RCs0kMQR1t7h RR=>"FGMs
";R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0FRmXh)bRFC0sNH
FM
-RR-8RQ:3Rp4
6RRkRVMHO0F"MRN"M8RR5p:QRAa);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0shRq7bRFC0sNH
FM
-RR-8RQ:3Rp4
nRRkRVMHO0F"MRN"M8RR5p:hRz1hQt R7;)RR:A2QaR0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDshRq7bRFC0sNH
FM
-RR-8RQ:3Rp4
(RRkRVMHO0F"MRFRs"5:pRRaAQ;RR):hRz1hQt R72skC0szMRht1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FRRm)FsbCNF0HMR

RR--QR8:pU34RR
RVOkM0MHFRs"F"pR5Rz:Rht1Qh; 7R:)RRaAQ2CRs0MksR1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNmsR)bRFC0sNH
FM
-RR-8RQ:3Rp4
gRRkRVMHO0F"MRM8NM"pR5RA:RQRa;)RR:zQh1t7h 2CRs0MksR1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFhsRqRh7FsbCNF0HMR

RR--QR8:pj3.RR
RVOkM0MHFRN"MMR8"5:pRR1zhQ th7);RRA:RQRa2skC0szMRht1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNRhhq7bRFC0sNH
FM
-RR-8RQ:3Rp.
4RRkRVMHO0F"MRM"FsRR5p:QRAa);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0smRh)bRFC0sNH
FM
-RR-8RQ:3Rp.
.RRkRVMHO0F"MRM"FsRR5p:hRz1hQt R7;)RR:A2QaR0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDsmRh)bRFC0sNH
FM
-RR-8RQ:3Rp.
dRRkRVMHO0F"MRG"FsRR5p:QRAa);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0smRX)bRFC0sNH
FM
-RR-8RQ:3Rp.
cRRkRVMHO0F"MRG"FsRR5p:hRz1hQt R7;)RR:A2QaR0sCkRsMzQh1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDsmRX)bRFC0sNH
FM
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3Rp.H6R#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3R.6
VRRk0MOHRFM"FGMs5"RpRR:A;QaR:)RR1zhQ th7s2RCs0kMhRz1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFsX)hmRCFbsHN0F
M
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR.p3n#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3Rp.
nRRkRVMHO0F"MRGsMF"pR5Rz:Rht1Qh; 7R:)RRaAQ2CRs0MksR1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNXsRhRm)FsbCNF0HMR

RR--QR8:p(3.RR
RVOkM0MHFRM"N85"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFsqRh7FsbCNF0HMR

RR--QR8:pU3.RR
RVOkM0MHFRM"N85"RpRR:1hQt R7;)RR:A2QaR0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNsqRh7FsbCNF0HMR

RR--QR8:pg3.RR
RVOkM0MHFRs"F"pR5RA:RQRa;)RR:1hQt R72skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFmsR)bRFC0sNH
FM
-RR-8RQ:3Rpd
jRRkRVMHO0F"MRFRs"5:pRRt1Qh; 7R:)RRaAQ2CRs0MksRt1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNRRm)FsbCNF0HMR

RR--QR8:p43dRR
RVOkM0MHFRN"MMR8"5:pRRaAQ;RR):QR1t7h 2CRs0MksRt1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FRhhq7bRFC0sNH
FM
-RR-8RQ:3Rpd
.RRkRVMHO0F"MRM8NM"pR5R1:RQ th7);RRA:RQRa2skC0s1MRQ th7R;
RR--)kC#D#0Rk$L0bRC:1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNhsRqRh7FsbCNF0HMR

RR--QR8:pd3dRR
RVOkM0MHFRF"Ms5"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFshRm)FsbCNF0HMR

RR--QR8:pc3dRR
RVOkM0MHFRF"Ms5"RpRR:1hQt R7;)RR:A2QaR0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNshRm)FsbCNF0HMR

RR--QR8:p63dRR
RVOkM0MHFRF"Gs5"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFsXRm)FsbCNF0HMR

RR--QR8:pn3dRR
RVOkM0MHFRF"Gs5"RpRR:1hQt R7;)RR:A2QaR0sCkRsM1hQt 
7;R-R-R#)CkRD0#0kL$:bCRt1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNsXRm)FsbCNF0HMR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp(3dRRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rdp3(RR
RMVkOF0HMGR"M"FsRR5p:QRAa);RR1:RQ th7s2RCs0kMQR1t7h ;R
R-)-RCD#k0kR#Lb0$C1:RQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0shRXmF)RbNCs0MHF
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RdUHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:pU3dRR
RVOkM0MHFRM"GFRs"5:pRRt1Qh; 7R:)RRaAQ2CRs0MksRt1Qh; 7
-RR-CR)#0kDRL#k0C$b:QR1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNRmXh)bRFC0sNH
FM
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpdHgR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
dgRkRVMHO0F"MRN"M8RR5p:QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa3
-RR-CR)#0kD:CR)#0kDRRFVN'M8HRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHjR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cjRkRVMHO0F"MRM8NM"pR5R1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A3QaRR
R-)-RCD#k0):RCD#k0VRFRMMN8M'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp43cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp34R
RVOkM0MHFRs"F"pR5R1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A3QaRR
R-)-RCD#k0):RCD#k0VRFR'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcH.R#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
c.RkRVMHO0F"MRM"FsRR5p:QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa3
-RR-CR)#0kD:CR)#0kDRRFVM'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHdR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cdRkRVMHO0F"MRG"FsRR5p:QR1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa3
-RR-CR)#0kD:CR)#0kDRRFVG'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHcR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
ccRkRVMHO0F"MRGsMF"pR5R1:RQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A3QaRR
R-)-RCD#k0):RCD#k0VRFRFGMsM'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp63cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp36R
RVOkM0MHFRM"N85"RpRR:zQh1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa3
-RR-CR)#0kD:CR)#0kDRRFVN'M8HRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHnR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cnRkRVMHO0F"MRM8NM"pR5Rz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAa
3RR-R-R#)Ck:D0R#)CkRD0FMVRN'M8HRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcH(R#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
c(RkRVMHO0F"MRFRs"5:pRR1zhQ th7s2RCs0kMQRAaR;
RR--)kC#D#0Rk$L0bRC:A3QaRR
R-)-RCD#k0):RCD#k0VRFR'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHUR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cURkRVMHO0F"MRM"FsRR5p:hRz1hQt R72skC0sAMRQ
a;R-R-R#)CkRD0#0kL$:bCRaAQ3RR
RR--)kC#DR0:)kC#DF0RVFRMsM'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpg3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3gR
RVOkM0MHFRF"Gs5"RpRR:zQh1t7h 2CRs0MksRaAQ;R
R-)-RCD#k0kR#Lb0$CA:RQRa3
-RR-CR)#0kD:CR)#0kDRRFVG'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3Rp6HjR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
6jRkRVMHO0F"MRGsMF"pR5Rz:Rht1Qh2 7R0sCkRsMA;Qa
-RR-CR)#0kDRL#k0C$b:QRAa
3RR-R-R#)Ck:D0R#)CkRD0FGVRM'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3

-RR-============================================================================R
R- -R8RoC7CC0OF0HMkRwMHO0F
M#R-R-============================================================================
R
R-Q-R8 :R3R4
RMVkOF0HMQR)1tQh_t 7 #R5HNoMD:R1RaAQ2CRs0MksRmAmph qRR=>"#sHC
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:CR)0Mks#)RazH RVMRNRCCPMH0R#CR800COCF8RMHR#oDMNRN1RM08RERC
RR--RRRRRRRRPkNDCERONCMo8sRVFNlRR''jRR0FN4R''
3
R-R-R:Q8R. 3
VRRk0MOHRFMwpqpQ_ht  7tRH5#oDMNRR1:A2QaR0sCkRsMApmm Rqh=">RVDND"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0R0)Ck#sMRza) VRHRRNMCMPC0#RHR08CCCO08MRFRo#HMRND1MRN8ER0CR
R-R-RRRRRRPRRNCDkRNOEM8oCRFVslRRN'R4'0NFRR''j3R

R-RR-============================================================================R
R-#-R0MsHoFROMsPC#MHFR8NMRHIs0FCRbNCs0MHF#R
R-=-==========================================================================R=
RR--0RECVDFDFMIHobRFC0sNH#FMRCNsRCbs8HCVM
C8RzRwhQBam0hRF0_#soHMRP5RNCDkRz:Rht1QhR 72 R)ahz)Rs#0H;Mo
wRRzahBQRmh0#F_0MsHoRR5PkNDCRR:1hQt R7RR)2R )azh0R#soHM;R

RR--CDGbH0OHD8$RCMVHCF8RbNCs0MHF#R

RHNDN0#RF#_L0MsHo#RHR_0F#H0sMroRzQh1t7h R0sCkRsM1Qa)h;t9
NRRD#HNR_0FLs#0HRMoH0#RF0_#soHMRQr1t7h R0sCkRsM1Qa)h;t9
NRRD#HNR_0FLNHMs#$_0MsHo#RHR_0F#H0sMroRzQh1t7h R0sCkRsM1Qa)h;t9
NRRD#HNR_0FLNHMs#$_0MsHo#RHR_0F#H0sMroR1hQt s7RCs0kMaR1)tQh9
;
RkRVMHO0F0MRF#_F0MsHoPR5NCDkRz:Rht1Qh2 7R0sCkRsM1Qa)h
t;RkRVMHO0F0MRF#_F0MsHoPR5NCDkR1:RQ th7s2RCs0kMaR1)tQh;R
RNNDH#FR0_0FON#D_0MsHo#RHR_0FFs#0HRMor1zhQ th7CRs0MksR)1aQ9ht;R
RNNDH#FR0_0FON#D_0MsHo#RHR_0FFs#0HRMort1QhR 7skC0s1MRah)Qt
9;
VRRk0MOHRFM0EF_#H0sM5oRPkNDCRR:zQh1t7h 2CRs0MksR)1aQ;ht
VRRk0MOHRFM0EF_#H0sM5oRPkNDCRR:1hQt R72skC0s1MRah)QtR;
RHNDN0#RFC_EG0_#soHMRRH#0EF_#H0sMroRzQh1t7h R0sCkRsM1Qa)h;t9
NRRD#HNR_0FE_CG#H0sMHoR#FR0_0E#soHMRQr1t7h R0sCkRsM1Qa)h;t9

RRCRM8h zv)_QBA;Qa
-
-=============================================================================-=
-=======================ROuN	CNoR8AF$=R======================================
==-=-=============================================================================

---B-RFsb$H0oER4�RgRg(LQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(dn3-g4g(-,
- RQ 1 R08NMNRs8ep]7RM1$0#ECHu#RNNO	o3C#RHaE#FR#kCsORDVHCNRl$FRM0CRL
R--OHFbCR8,#8FD,sRFROHMDCk88HRI0#ERFIV0NRsC00ENRRH##8FDR0IHE0FkRHIs0M0CR-
-RsbCl#H#HRFMVlsFRC0ER Q  0R1NNM8sR8#7NCbsC0lMR03a#EHRk#FsROCVCHDR$lN
R--LkCR#RC80HFRlCbDl0CMRH0E#0R#NNM8sN8RMl8RNL$RCHR8#H0sLCk08MRHRlOFbCHD8-
-RsVFlMRHR$NMRMlNMRCs#DFRFRMoN0#REOCRFHlbDRC8VlFsRC8F#FRM0DRNDRFI8CHsO-0
-CR8ObFlH0DNHRFMF0VREFCRsHHoMRND#sFkOVCRH3DCRHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--a#EHRObN	CNoR$lNRRLClHF8V8HCRR0FHDMOkR8CNH880MHFN8DRNR0NskCJH8sCRRL$0DFF#-,
-kRL00RHR#lk0MRHRRMFIRN$OMENo0CRECCRGs0CMRNDHCM0sOVNCF#RsHR#lNkD0MHFRELCNFPHs-
-RRFV0REC8OC#s0HbH3FMRRQ0Hb#RCHsl#L#HD0CRF8RN8FROlMlC0N#RMF8/s0RN0LsHk#0CR
0F-0-REbCRNNO	o8CRCNODsHN0F,M#R0LkR0MFRR0FOMENoFCRsCR8DCC0R$NMRHFsoNHMDHRDMRC#F-V
-ER0CNRbOo	NCCR8OsDNNF0HMa3REbCRNNO	oLCRFR8$lRN$LOCREoNMCF8RMRD$HNMROsOF8ONMC-
-R0IHEER0CCR0sRl#F(VR3N4RM(8R3F.RVER0H##R08NMN3s8

--b	NONRoCL$F8Rvhz B)Q_aAQR
H#
RRRR-R-R========================F=pORND1bkLssFoNRl#=================================R

RR--MDkDRMsNoNCRs$sNRMOF#M0N0
#
RFROMN#0Mh0Rq:zRR1zhQ th7R5j8MFI04FR2=R:R05FE#CsRR=>'2j';R
RO#FM00NMR1hqR1:RQ th7R5j8MFI04FR2RRR:5=RFC0Es=#R>jR''
2;
-RR-lRHblDCCNM00MHFRMOF0DsF#R

RMOF#M0N0mRh_)WqhtQhRA:Rm mpq:hR=NRVD;#CR-R-RV8CN0kDRR0FC0lHRsINMoHM#R

RMVkOF0HMQR1t7h _vhz_aAQ1qR5):tRRaQh )t 2CRs0MksRahqzp)qR
H#RRRRPHNsNCLDRQhAa:1RRahqzp)q;R
RRNRPsLHNDhCRRRRRRh:Rq)azq
p;RCRLo
HMRRRRHqVR)>tR=RRj0MEC
RRRRhRRRR:=q;)t
RRRR#CDCR
RRRRRh=R:Rq-5)4t+2R;
RCRRMH8RVR;
RhRRA1QaRR:=4R;
RIRRECHDR>hRRDjRF
FbRRRRRARhQRa1:h=RA1Qa+
4;RRRRRRRh:h=RR./R;R
RRMRC8FRDF
b;RRRRskC0shMRA1Qa;R
RCRM8VOkM0MHFRt1Qh_ 7h_zvA1Qa;R

RMVkOF0HMhRz1hQt h7_zAv_QRa15tq)Rh:Rq)azqRp2skC0shMRq)azqHpR#R
RRNRPsLHNDhCRA1QaRh:Rq)azq
p;RRRRPHNsNCLDRRhRR:RRRahqzp)q;R
RLHCoMR
RRRRh:q=R)
t;RRRRhaAQ1=R:R
4;RRRRIDEHCRRh>RR4DbFF
RRRRhRRA1QaRR:=haAQ1;+4
RRRRhRRRR:=hRR/.R;
RCRRMD8RF;Fb
RRRR0sCkRsMhaAQ1R;
R8CMRMVkOF0HMhRz1hQt h7_zAv_Q;a1
R
R-----------------------------------------------------------------------------R-
RR--0#EHR0HMCNsMDkRVMHO0FOMRFklb0RC#0RECNH880MHFRRFV0RIFzQh1t7h 
-RR-HRI0HERM0bkRsONsR$
RR--*ER0CIR0FsRNoCklMR0#NRsCF0VRE#CRNRlCDoCM0
E
RkRVMHO0FqMR7z7_ht1QhR 75Rp,)RR:zQh1t7h ;RRB:QRAas2RCs0kMhRz1hQt H7R#R
RRFROMN#0Mp0R_wp aRR:Q hatR ):p=R'MDCo-0E4R;
RNRRD#HNRRXpRRRRR:RRR1zhQ th7_5ppa wRI8FMR0FjH2R#;Rp
RRRRHNDNX#R)RRRRRRRRz:Rht1Qh5 7p _pw8aRF0IMF2RjRRH#)R;
RPRRNNsHLRDC)z 1p:aRR1zhQ th7_5ppa wRI8FMR0Fj
2;RRRRPHNsNCLDRQBAaRRR:QRAaRRRR=R:R
B;RCRLo
HMRRRRVRFsQMRHR0jRF_Rppa wRFDFbR
RRRRR)z 1pQa52=R:RQBAaFRGspRX5RQ2GRFsXQ)52R;
RRRRRQBAaRRRR:RR=BR5ARQaNRM8XQp52F2RsBR5ARQaNRM8XQ)52F2RsXR5p25QR8NMR5X)Q;22
RRRR8CMRFDFbR;
RsRRCs0kM R)1azp;R
RCRM8VOkM0MHFR7q7_1zhQ th7
;
R-R-RH0E#MRH0MCsNVDRk0MOHRFMObFlk#0CRC0ER8N8HF0HMVRFRF0IRt1Qh
 7R-R-R0IHEMRHbRk0OsNs$R
R-*-RRC0ERF0IRoNskMlC0N#RsFCRVER0CNR#lDCRC0MoER

RMVkOF0HM7Rq7Q_1t7h R,5pR:)RRt1Qh; 7R:BRRaAQ2CRs0MksRt1QhR 7HR#
RORRF0M#NRM0p _pw:aRRaQh )t RR:=pC'DMEo0-
4;RRRRNNDH#pRXRRRRRRRR:QR1t7h 5pp_ Rwa8MFI0jFR2#RHR
p;RRRRNNDH#)RXRRRRRRRR:QR1t7h 5pp_ Rwa8MFI0jFR2#RHR
);RRRRPHNsNCLDR1) zRpa:QR1t7h 5pp_ Rwa8MFI0jFR2R;
RPRRNNsHLRDCBaAQR:RRRaAQRRRRRR:=BR;
RoLCHRM
RVRRFQsRRRHMjFR0Rpp_ RwaDbFF
RRRR)RR p1za25QRR:=BaAQRsGFR5XpQG2RFXsR)25Q;R
RRRRRBaAQRRRRR=R:RA5BQNaRMX8Rp25Q2sRFRA5BQNaRMX8R)25Q2sRFRp5X5RQ2NRM8XQ)52
2;RRRRCRM8DbFF;R
RRCRs0MksR1) z;pa
CRRMV8Rk0MOHRFMq_771hQt 
7;
-RR-----------------------------------------------------------------------------R

RR--0#EHR0HMCNsMDsRbF8OCkRsCObFlk#0CR1zhQ th7HR8PHH#FRM
RR--oHHPM0oREJCRkHF0CRM0NRM8sNClHCM8sR3
RFbsOkC8s7CRQmev7hR5zRv,Xh7 m:vRR1zhQ th7X;RTazm,)RX QvqhRR:FRk0zQh1t7h 2#RH
RRRRsPNHDNLC RavRuRRz:Rht1Qh5 7h'zvDoCM08ERF0IMF2Rj;R
RRNRPsLHNDTCRzRmaRRR:zQh1t7h 5XvqQvvz5vhz'MDCo,0ER X7h'mvDoCM0-E24FR8IFM0R;j2
RRRRHNDN7#R vhmRRRRRz:Rht1Qh5 7Xh7 mDv'C0MoER-48MFI0jFR2#RHR X7h;mv
RRRRsPNHDNLCmRauaAQRQ:Rhta  
);RCRLo
HMRRRRau vR:RR=jR""z&hvR;
RTRRzRmaR=R:R05FE#CsRR=>'2j';R
RRmRauaAQRR:=-
4;RRRRVRFsKMRHRh7 msv'NCMoRFDFbR
RRRRRH7VR vhm5RK2=4R''ER0CRM
RRRRRaRRmQuAa=R:R
K;RRRRRRRRC0GH;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RR#RN#0CsRuamARQa>j=RRbsCFRs0"vhz B)Q_aAQ3e7Qv:m7Re7Q,mRv7F,Rs R)v$RLRsxCFR"
RRRRRP#CC0sH$sRCs;Fs
R
RRFRVsRRKHhMRzDv'C0MoEa-5mQuAa2+4RI8FMR0FjFRDFRb
RRRRRRHVau v5uamA+QaKR+48MFI0KFR2=R>R""j&h7 mav5mQuAaFR8IFM0RRj20MEC
RRRRRRRRva um5auaAQ+4K+RI8FMR0FK:2R=aR5 5vuaAmuQKa++84RF0IMF2RK2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR5""j&h7 mav5mQuAaFR8IFM0R2j2;R
RRRRRRzRTmKa52=R:R''4;R
RRRRRCRM8H
V;RRRRR#RN#0CsRva um5auaAQ+4K+2RR='
j'RRRRRRRRsFCbs"0Rh zv)_QBA3Qa7vQemR7:HCM0sDMNRsCsFHsRMER0CHR8PHH#FNMRDsoFHl0E"R
RRRRRRCR#PHCs0C$RsssF;R
RRMRC8FRDF
b;RRRRXmTzaRRR:)=R Z1Q z5TmRa,XmTzaC'DMEo02R;
RXRR)q vQ:hR= R)1 QZ5va uX,R)q vQDh'C0MoE
2;RMRC8sRbF8OCkRsC7vQem
7;
-RR----------------pNFODkR1LFbsolsN#RR-#VEH0F/s0CN0R#Fb-------------------------R

RMVkOF0HM1RXp5pRqR)t:QRAa _eB)am;mRBzRha:qRhaqz)ps2RCs0kMQRAa _eB)amR
H#RRRRO#FM00NMRtq)_RpR:hRQa  t)RRRRRRRRRRRRRRRRRRRRR:=q')tDoCM04E-;R
RRDRNHRN#Xtq)RRRRRRR:A_Qaea Bmq)5)pt_RI8FMR0FjH2R#)RqtR;
RPRRNNsHLRDC)z 1p:aRRaAQ_Be a5m)q_)tpFR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRHBVRmazhRR<=q_)tpER0CRM
RRRRR1) z5paq_)tpFR8IFM0RzBmhRa2:X=Rq5)tq_)tpm-BzRha8MFI0jFR2R;
RCRRMH8RVR;
RsRRCs0kM R)1azp;R
RCRM8VOkM0MHFRpX1p
;
RkRVMHO0FXMR1R)p5tq)RA:RQea_ mBa)B;RmazhRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
RRRRMOF#M0N0)RqtR_pRQ:Rhta  R)RRRRRRRRRRRRRRRRRR=R:Rtq)'MDCo-0E4R;
RNRRD#HNR)XqtRRRR:RRRaAQ_Be a5m)q_)tpFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDR1) zRpa:QRAa _eB)am5tq)_8pRF0IMF2RjRR:=5EF0CRs#='>Rj;'2
LRRCMoH
RRRRRHVBhmza=R<Rtq)_0pRE
CMRRRRR R)1azp5tq)_Bp-mazhRI8FMR0Fj:2R=qRX)qt5)pt_RI8FMR0FBhmza
2;RRRRCRM8H
V;RRRRskC0s)MR p1zaR;
R8CMRMVkOF0HM1RX)
p;
VRRk0MOHRFMXq1)R)5qtRR:A_Qaea BmR);BhmzaRR:hzqa)2qpR0sCkRsMA_Qaea BmH)R#R
RRFROMN#0Mq0R)pt_RRR:Q hatR ):q=R)Dt'C0MoE;-4
RRRRHNDNX#RqR)tRRRRRA:RQea_ mBa))5qtR_p8MFI0jFR2#RHRtq);R
RRNRPsLHND)CR p1zaRR:A_Qaea Bmq)5)pt_RI8FMR0Fj
2;RRRRPHNsNCLDRmXBzRha:qRhaqz)p=R:RzBmh
a;RCRLo
HMRRRRH5VR5tq)'MDCoR0E<4=R2sRFRB5XmazhRj=R202RERCMskC0sqMR)
t;RRRRCCD#
RRRRHRRVXR5BhmzaRR>q_)tp02RERCMXzBmhRaRRRRRRRRRRR:=q_)tpR;
RRRRR8CMR;HV
RRRR)RR p1za)5qt-_pXzBmh8aRF0IMF2RjRRRRRRRRRRRRRR:=Xtq)5tq)_8pRF0IMFBRXmazh2R;
RRRRR1) z5paq_)tpFR8IFM0R)5qtR_p-BRXmazhR4+R2:2R=FR50sEC#>R=R)Xqt)5qt2_p2R;
RCRRMH8RVR;
RsRRCs0kM R)1azp;R
RCRM8VOkM0MHFR)X1q
;
RkRVMHO0FXMR)Rmp5tq)RA:RQea_ mBa)B;RmazhRh:Rq)azqRp2skC0sAMRQea_ mBa)#RH
RRRRMOF#M0N0)RqtR_pRQ:Rhta  R)RRRRRRRRRRRRRRRRRR=R:Rtq)'MDCo-0E4R;
RNRRD#HNR)XqtRRRR:RRRaAQ_Be a5m)q_)tpFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDR1) zRpa:QRAa _eB)am5tq)_8pRF0IMF2RjRR:=Xtq);R
RRNRPsLHNDBCRmazhvRR:Q hat; )
LRRCMoH
RRRRzBmhRav:B=RmazhR8lFR)5qtR_p+2R4;R
RRVRHRzBmhRav/j=RRC0EMR
RRRRR)z 1pqa5)pt_RI8FMR0FBhmzaRv2:X=Rq5)tq_)tpm-BzvhaRI8FMR0Fj
2;RRRRR R)1azp5zBmh-av4FR8IFM0RRj2R=R:R)Xqt)5qtR_p8MFI0qFR)pt_-zBmh+av4
2;RRRRCRM8H
V;RRRRskC0s)MR p1zaR;
R8CMRMVkOF0HM)RXm
p;
VRRk0MOHRFMX))mR)5qtRR:A_Qaea BmR);BhmzaRR:hzqa)2qpR0sCkRsMA_Qaea BmH)R#R
RRFROMN#0Mq0R)pt_RRR:Q hatR )RRRRRRRRRRRRRRRRR:RR=)RqtC'DMEo0-
4;RRRRNNDH#qRX)RtRRRRR:QRAa _eB)am5tq)_8pRF0IMF2RjRRH#q;)t
RRRRsPNHDNLC R)1azpRA:RQea_ mBa))5qtR_p8MFI0jFR2=R:R)XqtR;
RPRRNNsHLRDCBhmza:vRRaQh )t ;R
RLHCoMR
RRmRBzvhaRR:=BhmzaFRl8qR5)pt_R4+R2R;
RHRRVmRBzvhaRR/=jER0CRM
RRRRR1) z5paq_)tpm-BzvhaRI8FMR0FjR2RRRRRRR:=Xtq)5tq)_8pRF0IMFmRBzvha2R;
RRRRR1) z5paq_)tpFR8IFM0Rtq)_Bp-mazhv2+4RR:=Xtq)5zBmh-av4FR8IFM0R;j2
RRRR8CMR;HV
RRRR0sCkRsM)z 1p
a;RMRC8kRVMHO0FXMR);m)
R
R----------------ROpFN1DRksLbFNosl-#RRD)CNF0HMRNDmsbCNs0F#-R------------------
-
R-R-
-RR-CRtMNCsD=R""FRVshRz1hQt P7RCFO0sR#,#CNlRMDCo
0ER-R-
VRRk0MOHRFMzQh1t7h _z Tq5pRp),RRz:Rht1Qh2 7R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMQRAa _eB)am5Rp2=QRAa _eB)am5;)2
CRRMV8Rk0MOHRFMzQh1t7h _z Tq
p;
-RR-R
R-t-RCsMCN"DR=V"RF1sRQ th7CRPOs0F##,RNRlCDoCM0RE
R
--RkRVMHO0F1MRQ th7T_ zRqp5Rp,)RR:1hQt R72skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRaAQ_Be a5m)p=2RRaAQ_Be a5m))
2;RMRC8kRVMHO0F1MRQ th7T_ z;qp
R
R-R-
RR--tCCMsRND"R<"VRFszQh1t7h ROPC0#Fs,NR#lDCRC0MoER
R-R-
RMVkOF0HMhRz1hQt p7_ R115Rp,)RR:zQh1t7h 2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0sAMRQea_ mBa)25pRA<RQea_ mBa)25);R
RCRM8VOkM0MHFR1zhQ th7 _p1
1;
-RR-R
R-t-RCsMCN"DR<V"Rk0MOHRFMVRFs1hQt P7RCFO0sR#,#CNlRMDCo
0ER-R-
VRRk0MOHRFM1hQt p7_ R115Rp,)RR:1hQt R72skC0sAMRm mpqHhR#R
RR-R-RChC8DRNHCN##FR0R#N#kRsCHCM8GHR8s0COH
FMRRRRPHNsNCLDRaQh _)hpRR:1hQt j75RR0FpC'DMEo0-;42
RRRRsPNHDNLChRQah )_:)RRt1Qh5 7jFR0RD)'C0MoE2-4;R
RLHCoMR
RRhRQah )_RpRR=R:R
p;RRRRQ ha))h_RRRR:)=R;R
RRhRQah )_jp52=R:R0MFRaQh _)hp25j;R
RRhRQah )_j)52=R:R0MFRaQh _)h)25j;R
RRCRs0MksRaAQ_Be a5m)Q ha)ph_2RR<A_Qaea BmQ)5h)a h2_);R
RCRM8VOkM0MHFRt1Qh_ 7p1 1;R

R
--R-R-RMtCCDsNR="<"kRVMHO0FVMRFzsRht1QhR 7P0COF,s#Rl#NCCRDMEo0
-RR-R
RVOkM0MHFR1zhQ th7 _p1m1_)T_ zRqp5Rp,)RR:zQh1t7h 2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0sAMRQea_ mBa)25pRR<=A_Qaea Bm))52R;
R8CMRMVkOF0HMhRz1hQt p7_ _11m )_Tpzq;R

R
--R-R-RMtCCDsNR="<"kRVMHO0FVMRF1sRQ th7CRPOs0F##,RNRlCDoCM0RE
R
--RkRVMHO0F1MRQ th7 _p1m1_)T_ zRqp5Rp,)RR:1hQt R72skC0sAMRm mpqHhR#R
RR-R-RChC8DRNHCN##FR0R#N#kRsCHCM8GHR8s0COH
FMRRRRPHNsNCLDRaQh _)hpRR:1hQt j75RR0FpC'DMEo0-;42
RRRRsPNHDNLChRQah )_:)RRt1Qh5 7jFR0RD)'C0MoE2-4;R
RLHCoMR
RRhRQah )_RpRRRRRRRRRRRRRRRRRR=R:R
p;RRRRQ ha))h_RRRRRRRRRRRRRRRRRRRR:)=R;R
RRhRQah )_jp52RRRRRRRRRRRRRRRR=R:R0MFRaQh _)hp25j;R
RRhRQah )_j)52RRRRRRRRRRRRRRRR=R:R0MFRaQh _)h)25j;R
RRCRs0MksRaAQ_Be a5m)Q ha)ph_2=R<RaAQ_Be a5m)Q ha))h_2R;
R8CMRMVkOF0HMQR1t7h _1p 1)_m_z Tq
p;
V
Sk0MOHRFMMLklCFs_VH_L0k#_Mo#HM5C8MRkl:NRM0NksDs2RCs0kMNRM0NksD#RH
PSSNNsHLRDC0,lbRlMkL_CsFLV_HR0#:NRM0NksDS;
LHCoMS
S0Rlb:M=Rk
l;SkSMlsLC__FVL#H0RR:=4S;
SHIED0CRl>bRRD4RF
FbSMSSkClLsV_F_0LH#=R:RlMkL_CsFLV_H+0#4S;
SlS0b=R:Rb0l/
.;SMSC8FRDF
b;SCSs0MksRlMkL_CsFLV_H;0#
MSC8kRMlsLC__FVL#H0_#kMHCoM8S;
VOkM0MHFRlMkL_CsFLV_H_0##MHoC58RM:klR0HMCsoC2CRs0MksR0MNkDsNR
H#SNSPsLHNDMCRkClLsV_F_0LH#M:RNs0kN
D;SNSPsLHND0CRlRb:MkN0s;ND
CSLo
HMSlS0b=R:RlMk;S
SHMVRk<lRR0jRE
CMSRSR0Rlb:-=R5lMk+;42
CSSMH8RVS;
SlMkL_CsFLV_HR0#:4=R;S
SIDEHClR0bRR>jFRDFSb
SMRRkClLsV_F_0LH#=R:RlMkL_CsFLV_H+0#4S;
S0RRl:bR=lR0bRR/.S;
S8CMRFDFbS;
S0sCkRsMMLklCFs_VH_L0
#;S8CMRlMkL_CsFLV_H_0##MHoC
8;
RRR-=-R=====================GR b0FsCw8Rk0MOH#FMR================================
==
RRRRMVkOF0HMqR"A51"p1:RQ th7s2RCs0kMQR1t7h R
H#SNSPsLHNDsCRCD#k01:RQ th7'5pDoCM04E-RI8FMR0Fj
2;RRRRLHCoMS
SH5VRp'5pD0CV2RR='2j'RC0EMS
SS#sCkRD0:p=R;S
SCCD#
SSSskC#D:0R=jRRRp-R;S
SCRM8H
V;RRRRRRRRskC0ssMRCD#k0R;
RCRRM
8;
RRRRMVkOF0HMCRs#CHxR)5qt1:RQ th7h;R 1W_Q:Z Rahqzp)q2CRs0MksRt1QhR 7HR#
RRRRRRRRRNRRD#HNR0LH#1:RQ th7)5qt 'ph]ta-84RF0IMF2RjRRH#q;)t
RRRRRRRRRRRRsPNHDNLCCRs#0kD:QR1t7h 5Wh _Z1Q R-48MFI0jFR2=R:R05FE#CsRR=>'2j';R
RRRRRRRRRRFROMN#0MN0RsCopMQ:Rhta  :)R=)Rqt 'ph]ta;R
RRCRLo
HMRRRRRRRRRRRRH5VRNpsoC=MRRWh _Z1Q 02RE
CMRRRRRRRRRRRRRRRRR0sCkRsML#H0;R
RRRRRRRRRRMRC8VRH;R

RRRRRRRRRsRRCD#k0=R:R05FE#CsRR=>q5)tq')tpa w2
2;RRRRRRRRRRRRH5VRh_ W1 QZR.<RRRFsNpsoC<MRRR.20MEC
RRRRRRRRRRRRRRRR0sCkRsMskC#D
0;RRRRRRRRRRRRCHD#VNR5sCopMRR<h_ W1 QZ2ER0CRM
RRRRRRRRRRRRRRRRskC#DN05sCopMR-.8MFI0jFR2=R:R0LH#s5NoMpC-8.RF0IMF2Rj;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRRRRRskC#Dh05 1W_Q-Z .FR8IFM0RRj2:L=RH50#h_ W1 QZ-8.RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRRRRRCRs0MksR#sCk;D0
RRRR8CM;S

VOkM0MHFR""<R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMa )z;S
SCRM8H
V;SCSs0MksR""<5Rp,azm_ht1Qh5 7)p,R'hp t2a]2S;
C;M8
V
Sk0MOHRFM"R<"5Rp:hzqa);qpRR):zQh1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0k#_Mo#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0swMRq p1;S
SCRM8H
V;SCSs0MksR""<5_amzQh1t7h 5Rp,) 'ph]ta2),R2S;
C;M8
V
Sk0MOHRFM"R<"5Rp:Q hat; )RR):1hQt R72skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_o#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0spMRRj<R;S
SCRM8H
V;SCSs0MksR""<5_am1hQt p75,'R)pt ha,]2R;)2
MSC8<R""
;
SMVkOF0HM<R"":5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMjRR<)S;
S8CMR;HV
sSSCs0kM<R"",5pR_am1hQt )75,'Rppt ha2]2;C
SM"8R<
";
kSVMHO0F"MR<R="5Rp:zQh1t7h ;:R)Rahqzp)q2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0k#_Mo#HM5C8)
2;SVSHRlMkL#H0Rp>R'hp tRa]0MEC
SSSskC0saMR);z 
CSSMH8RVS;
S0sCkRsM""<=5Rp,azm_ht1Qh5 7)p,R'hp t2a]2S;
C;M8
V
Sk0MOHRFM""<=R:5pRahqzp)q;:R)R1zhQ th7s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;p2
HSSVkRMl0LH#RR>) 'ph]taRC0EMS
SS0sCkRsMw1qp S;
S8CMR;HV
sSSCs0kM<R"=a"5mh_z1hQt p75,'R)pt ha,]2R;)2
MSC8
;
SMVkOF0HM<R"=5"RpQ:Rhta  R);)1:RQ th7s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0##MHoCp852S;
SRHVMLklHR0#>'R)pt ha0]RE
CMSsSSCs0kMRRp<;Rj
CSSMH8RVS;
S0sCkRsM""<=5_am1hQt p75,'R)pt ha,]2R;)2
MSC8<R"=
";
kSVMHO0F"MR<5="p1:RQ th7);R:hRQa  t)s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0##MHoC)852S;
SRHVMLklHR0#>'Rppt ha0]RE
CMSsSSCs0kMRRj<;R)
CSSMH8RVS;
S0sCkRsM""<=5Rp,a1m_Q th7,5)Rpp' aht];22
MSC8<R"=
";
R
RRRRRVOkM0MHFR"">R:5pR1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMw1qp S;
S8CMR;HV
sSSCs0kM>R"",5pR_amzQh1t7h 5R),p 'ph]ta2
2;S8CM;S

VOkM0MHFR"">R:5pRahqzp)q;:R)R1zhQ th7s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;p2
HSSVkRMl0LH#RR>) 'ph]taRC0EMS
SS0sCkRsMa )z;S
SCRM8H
V;SCSs0MksR"">5_amzQh1t7h 5Rp,) 'ph]ta2),R2S;
C;M8
V
Sk0MOHRFM"R>"5Rp:Q hat; )RR):1hQt R72skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_o#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0spMRRj>R;S
SCRM8H
V;SCSs0MksR"">5_am1hQt p75,'R)pt ha,]2R;)2
MSC8>R""
;
SMVkOF0HM>R"":5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMjRR>)S;
S8CMR;HV
sSSCs0kM>R"",5pR_am1hQt )75,'Rppt ha2]2;C
SM"8R>
";
R
RRRRRVOkM0MHFR=">"pR5:hRz1hQt R7;)h:Rq)azqRp2skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_#kMHCoM825);S
SHMVRkHlL0>#RRpp' aht]ER0CSM
SCSs0MksRpwq1
 ;SMSC8VRH;S
SskC0s"MR>5="pa,Rmh_z1hQt )75,'Rppt ha2]2;C
SM
8;
kSVMHO0F"MR>R="5Rp:hzqa);qpRR):zQh1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0k#_Mo#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0saMR);z 
CSSMH8RVS;
S0sCkRsM"">=5_amzQh1t7h 5Rp,) 'ph]ta2),R2S;
C;M8
V
Sk0MOHRFM"">=R:5pRaQh )t ;:R)Rt1Qh2 7R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;p2
HSSVkRMl0LH#RR>) 'ph]taRC0EMS
SS0sCkRsMpRR>jS;
S8CMR;HV
sSSCs0kM>R"=a"5mQ_1t7h 5Rp,) 'ph]ta2),R2S;
CRM8"">=;S

VOkM0MHFR=">":5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMjRR>)S;
S8CMR;HV
sSSCs0kM>R"=p"5,mRa_t1Qh5 7)p,R'hp t2a]2S;
CRM8"">=;


SMVkOF0HM=R"":5pRt1Qh; 7RR):Q hat2 )R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;)2
HSSVk5Ml0LH#RR>p 'ph]ta2ER0CSM
SCSs0Mks5pwq1; 2
CSSD
#CSsSSCs0kM=R"",5pR_am1hQt )75,'Rppt ha2]2;S
SCRM8H
V;S8CMR""=;

SSMVkOF0HM=R"":5pRaQh )t ;:R)Rt1Qh2 7R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;p2
HSSVk5Ml0LH#RR>) 'ph]ta2ER0CSM
SCSs0Mks5pwq1; 2
CSSD
#CSsSSCs0kM=R"",5)R_am1hQt p75,'R)pt ha2]2;S
SCRM8H
V;S8CMR""=;R

RRRRRMVkOF0HM=R"":5pR1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;)2
HSSVk5Ml0LH#RR>p 'ph]ta2ER0CSM
SCSs0Mks5pwq1; 2
CSSD
#CSsSSCs0kM=R"",5pR_amzQh1t7h 5R),p 'ph]ta2
2;SMSC8VRH;C
SM"8R=
";SV
Sk0MOHRFM"5="ph:Rq)azqRp;)z:Rht1Qh2 7R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#M_k#MHoCp852S;
S5HVMLklHR0#>'R)pt haR]20MEC
SSSskC0swM5q p12S;
S#CDCS
SS0sCkRsM"5=")a,Rmh_z1hQt p75,'R)pt ha2]2;S
SCRM8H
V;S8CMR""=;

SSMVkOF0HMlR"FR8"5Rp,)1:RQ th7s2RCs0kMQR1t7h R
H#SsPNHDNLCCRs#0kDR#:RHCoM8'5)DoCM04E-RI8FMR0Fj
2;SsPNHDNLCCRslMNH8RCs:MRk#MHoC)85'MDCo-0E4FR8IFM0R;j2
NSPsLHND0CRlRbD:MRk#MHoCp85'MDCo-0E4FR8IFM0R;j2
NSPsLHND0CRlRbs:MRk#MHoC)85'MDCo-0E4FR8IFM0R;j2
NSPsLHNDICRHE80NRR:HCM0oRCs:p=R'MDCo;0E
NSPsLHNDICRHE80LRR:HCM0oRCs:)=R'MDCo;0E
NSPsLHNDsCRH0oEM:CoRmAmph qRR:=w1qp S;
LHCoMS
SH5VRp'5ppa w2RR='24'RC0EMS
SSb0lD=R:R#kMHCoM8p5-2S;
S#CDCS
SSb0lD=R:R#kMHCoM825p;S
SCRM8H
V;SVSHR55)) 'pwRa2=4R''02RE
CMS0SSlRbs:k=RMo#HM5C8-;)2
SSSsEHo0oMCRR:=a )z;S
SCCD#
SSS0slbRR:=kHM#o8MC5;)2
CSSMH8RVS;
S5HV)RR=j02RE
CMSsSSCD#k0=R:R05FE#CsRR=>'2j';S
SCCD#SSR
S-S-sNClHCM8sS
SSlsCN8HMC:sR=sR"C5l"0Dlb,b0ls
2;SHSSVHRsoME0CNoRMp8R5pp' 2wa=''4RC0EMS
SSsRRCHlNMs8CRR:="-j"sNClHCM8sS;
SDSC#RHVsEHo0oMCR8NMRlsCN8HMC=s/"Rj"0MEC
SSSRCRslMNH8RCs:s=RCHlNMs8C-b0lsS;
SDSC#RHVp'5ppa w24=''MRN8CRslMNH8/Cs=""jRC0EMS
SSsRRCHlNMs8CRR:=0slb-lsCN8HMC
s;SSSSCRM8H
V;SsSSCD#k0=R:Rt1Qh5 7sNClHCM8s
2;SMSC8VRH;S
SskC0ssMRCD#k0S;
CRM8"8lF"
;
RRRR-=-R=========================================================================
==R-R-R:Q8Rdq3gR
RVOkM0MHFRMVH8C_DVF0l#50RqR)t:hRz1hQt R7;YRR:A2QaR0sCkRsMQ hatR )HR#
RoLCHRM
RVRRFQsRhX7 RRHMq')tsoNMCFRDFRb
RRRRRRHVq5)tQ h7X=2RR0YRE
CMRRRRRRRRskC0sQMRhX7 ;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RRCRs0MksR;-4
CRRMV8Rk0MOHRFMV8HM_VDC0#lF0
;
R-R-R:Q8Rcq3jR
RVOkM0MHFRMVH8C_DVF0l#50RqR)t:QR1t7h ;RRY:QRAas2RCs0kMhRQa  t)#RH
LRRCMoH
RRRRsVFR7Qh HXRM)RqtN'sMRoCDbFF
RRRRHRRV)Rqth5Q72 XRY=RRC0EMR
RRRRRRCRs0MksR7Qh 
X;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRRskC0s-MR4R;
R8CMRMVkOF0HMHRVMD8_ClV0F;#0
R
R-Q-R8q:R3
c4RkRVMHO0FVMRH_M8sEHo0#lF0qR5):tRR1zhQ th7Y;RRA:RQRa2skC0sQMRhta  H)R#R
RLHCoMR
RRFRVshRQ7R XHqMR)st'CsPC#sC_NCMoRFDFbR
RRRRRHqVR)Qt5hX7 2RR=YER0CRM
RRRRRsRRCs0kMhRQ7; X
RRRRCRRMH8RVR;
RCRRMD8RF;Fb
RRRR0sCkRsM-
4;RMRC8kRVMHO0FVMRH_M8sEHo0#lF0
;
R-R-R:Q8Rcq3.R
RVOkM0MHFRMVH8H_solE0FR#05tq)R1:RQ th7Y;RRA:RQRa2skC0sQMRhta  H)R#R
RLHCoMR
RRFRVshRQ7R XHqMR)st'CsPC#sC_NCMoRFDFbR
RRRRRHqVR)Qt5hX7 2RR=YER0CRM
RRRRRsRRCs0kMhRQ7; X
RRRRCRRMH8RVR;
RCRRMD8RF;Fb
RRRR0sCkRsM-
4;RMRC8kRVMHO0FVMRH_M8sEHo0#lF0
;
R-R-R:Q8RdB3(R
RVOkM0MHFRhvQQvvzR,5pR:)RR1zhQ th7s2RCs0kMhRz1hQt H7R#R
RRFROMN#0M10RQRZ :qRhaqz)p=R:RXvqQvvz5Dp'C0MoE),R'MDCo20E;R
RLHCoMR
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MECR0sCkRsMh;qz
RRRR8CMR;HV
RRRRRHVzQh1t7h _1p 1 5)1 QZ5Rp,1 QZ2),R Z1Q ,5)RZ1Q R220MEC
RRRRsRRCs0kM R)1 QZ5Rp,1 QZ2R;
RCRRD
#CRRRRRCRs0MksR1) Q5Z )1,RQ2Z ;R
RRMRC8VRH;R
RCRM8VOkM0MHFRhvQQvvz;R

RR--QR8:BU3d
VRRk0MOHRFMvQQhvRzv5Rp,)RR:1hQt R72skC0s1MRQ th7#RH
RRRRMOF#M0N0QR1Z: RRahqzp)qRR:=vQqXv5zvpC'DMEo0,'R)DoCM0;E2
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RERCMskC0shMRq
1;RRRRCRM8H
V;RRRRH1VRQ th7 _p1)15 Z1Q ,5pRZ1Q R2,)Q 1Z) 5,QR1Z2 2RC0EMR
RRRRRskC0s)MR Z1Q ,5pRZ1Q 
2;RRRRCCD#
RRRRsRRCs0kM R)1 QZ5R),1 QZ2R;
RCRRMH8RVR;
R8CMRMVkOF0HMQRvhzQvv
;
R-R-R:Q8RdB3gR
RVOkM0MHFRhvQQvvzRR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h R
H#RCRLo
HMRRRRskC0svMRQvhQzav5mh_z1hQt p75,'R)DoCM0,E2R;)2
CRRMV8Rk0MOHRFMvQQhv;zv
R
R-Q-R8B:R3
cjRkRVMHO0FvMRQvhQz5vRpRR:Q hat; )R:)RRt1Qh2 7R0sCkRsM1hQt H7R#R
RLHCoMR
RRCRs0MksRhvQQvvz5_am1hQt p75,'R)DoCM0,E2R;)2
CRRMV8Rk0MOHRFMvQQhv;zv
R
R-Q-R8B:R3
c4RkRVMHO0FvMRQvhQz5vRpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMhRz1hQt H7R#R
RLHCoMR
RRCRs0MksRhvQQvvz5Rp,azm_ht1Qh5 7)p,R'MDCo20E2R;
R8CMRMVkOF0HMQRvhzQvv
;
R-R-R:Q8RcB3.R
RVOkM0MHFRhvQQvvzRR5p:QR1t7h ;RR):hRQa  t)s2RCs0kMQR1t7h R
H#RCRLo
HMRRRRskC0svMRQvhQzpv5,mRa_t1Qh5 7)p,R'MDCo20E2R;
R8CMRMVkOF0HMQRvhzQvv
;
R-R-R============================================================================R

RR--QR8:Bd3c
VRRk0MOHRFMvQqXvRzv5Rp,)RR:zQh1t7h 2CRs0MksR1zhQ th7#RH
RRRRMOF#M0N0QR1Z: RRahqzp)qRR:=vQqXv5zvpC'DMEo0,'R)DoCM0;E2
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RERCMskC0shMRq
z;RRRRCRM8H
V;RRRRHzVRht1Qh_ 7p1 151) Q5Z p1,RQ2Z , R)1 QZ5R),1 QZ202RE
CMRRRRRCRs0MksR1) Q5Z )1,RQ2Z ;R
RRDRC#RC
RRRRR0sCkRsM)Q 1Zp 5,QR1Z; 2
RRRR8CMR;HV
CRRMV8Rk0MOHRFMvQqXv;zv
R
R-Q-R8B:R3
ccRkRVMHO0FvMRqvXQz5vRp),RR1:RQ th7s2RCs0kMQR1t7h R
H#RRRRO#FM00NMRZ1Q RR:hzqa)Rqp:v=RqvXQzpv5'MDCo,0ERD)'C0MoE
2;RCRLo
HMRRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CsMRCs0kMqRh1R;
RCRRMH8RVR;
RHRRVQR1t7h _1p 1 5)1 QZ5Rp,1 QZ2),R Z1Q ,5)RZ1Q R220MEC
RRRRsRRCs0kM R)1 QZ5R),1 QZ2R;
RCRRD
#CRRRRRCRs0MksR1) Q5Z p1,RQ2Z ;R
RRMRC8VRH;R
RCRM8VOkM0MHFRXvqQvvz;R

RR--QR8:B63c
VRRk0MOHRFMvQqXvRzv5:pRRahqzp)q;RR):hRz1hQt R72skC0szMRht1QhR 7HR#
RoLCHRM
RsRRCs0kMqRvXzQvvm5a_1zhQ th7,5pRD)'C0MoER2,)
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcRn
RMVkOF0HMqRvXzQvvpR5RQ:Rhta  R);)RR:1hQt R72skC0s1MRQ th7#RH
LRRCMoH
RRRR0sCkRsMvQqXv5zva1m_Q th7,5pRD)'C0MoER2,)
2;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcR(
RMVkOF0HMqRvXzQvvpR5Rz:Rht1Qh; 7R:)RRahqzp)q2CRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMvQqXv5zvpa,Rmh_z1hQt )75,'RpDoCM02E2;R
RCRM8VOkM0MHFRXvqQvvz;R

RR--QR8:BU3c
VRRk0MOHRFMvQqXvRzv5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMqRvXzQvv,5pR_am1hQt )75,'RpDoCM02E2;R
RCRM8VOkM0MHFRXvqQvvz;R

RR--============================================================================
R
R-Q-R8B:R3
cgRkRVMHO0F"MR?R>"5Rp,)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRR)>RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R">
";
-RR-8RQ:3RB6Rj
RMVkOF0HM?R">5"Rp),RR1:RQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR>)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;>"
R
R-Q-R8B:R3
64RkRVMHO0F"MR?R>"5:pRRahqzp)q;RR):hRz1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRVRHR>pRR0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:B.36
VRRk0MOHRFM""?>RR5p:hRQa  t));RR1:RQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR>)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;>"
R
R-Q-R8B:R3
6dRkRVMHO0F"MR?R>"5:pRR1zhQ th7);RRh:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRVRHR>pRR0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:Bc36
VRRk0MOHRFM""?>RR5p:QR1t7h ;RR):hRQa  t)s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR>)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;>"
R
R-=-R=========================================================================
==
-RR-8RQ:3RB6R6
RMVkOF0HM?R"<5"Rp),RRz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RHRRVRRp<RR)0MEC
RRRRsRRCs0kM4R''R;
RCRRD
#CRRRRRCRs0MksR''j;R
RRMRC8VRH;R
RCRM8VOkM0MHFR<"?"
;
R-R-R:Q8R6B3nR
RVOkM0MHFR<"?"pR5,RR):QR1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRR)<RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
-RR-8RQ:3RB6R(
RMVkOF0HM?R"<5"RpRR:hzqa);qpR:)RR1zhQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR<)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
6URkRVMHO0F"MR?R<"5:pRRaQh )t ;RR):QR1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRR)<RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
-RR-8RQ:3RB6Rg
RMVkOF0HM?R"<5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR<)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
njRkRVMHO0F"MR?R<"5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRR)<RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
-RR-=R==========================================================================
=
R-R-R:Q8RnB34R
RVOkM0MHFR<"?=5"Rp),RRz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RHRRVRRp<)=RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
n.RkRVMHO0F"MR?"<=R,5pR:)RRt1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RHRRVRRp<)=RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
ndRkRVMHO0F"MR?"<=RR5p:qRhaqz)p);RRz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RHRRVRRp<)=RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
ncRkRVMHO0F"MR?"<=RR5p:hRQa  t));RR1:RQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVp=R<R0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?<"
;
R-R-R:Q8RnB36R
RVOkM0MHFR<"?=5"RpRR:zQh1t7h ;RR):qRhaqz)ps2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVp=R<R0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?<"
;
R-R-R:Q8RnB3nR
RVOkM0MHFR<"?=5"RpRR:1hQt R7;)RR:Q hat2 )R0sCkRsMARQaHR#
RoLCHRM
RHRRVRRp<)=RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
R-=-R=========================================================================
==
-RR-8RQ:3RBnR(
RMVkOF0HM?R">R="5Rp,)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR>=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?">=;R

RR--QR8:BU3n
VRRk0MOHRFM"=?>"pR5,RR):QR1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR>=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?">=;R

RR--QR8:Bg3n
VRRk0MOHRFM"=?>"pR5Rh:Rq)azqRp;)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR>=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?">=;R

RR--QR8:Bj3(
VRRk0MOHRFM"=?>"pR5RQ:Rhta  R);)RR:1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRVRHR>pR=RR)0MEC
RRRRsRRCs0kM4R''R;
RCRRD
#CRRRRRCRs0MksR''j;R
RRMRC8VRH;R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RB(R4
RMVkOF0HM?R">R="5:pRR1zhQ th7);RRh:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRVRHR>pR=RR)0MEC
RRRRsRRCs0kM4R''R;
RCRRD
#CRRRRRCRs0MksR''j;R
RRMRC8VRH;R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RB(R.
RMVkOF0HM?R">R="5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR>=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?">=;R

RR--============================================================================
R
R-Q-R8B:R3
(dRkRVMHO0F"MR?R="5Rp,)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRR)=RRC0EMR
RRRRRskC0s'MR4
';RRRRCCD#
RRRRsRRCs0kMjR''R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(Rc
RMVkOF0HM?R"=5"Rp),RR1:RQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;="
R
R-Q-R8B:R3
(6RkRVMHO0F"MR?R="5:pRRahqzp)q;RR):hRz1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRVRHR=pRR0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?=;R

RR--QR8:Bn3(
VRRk0MOHRFM""?=RR5p:hRQa  t));RR1:RQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;="
R
R-Q-R8B:R3
((RkRVMHO0F"MR?R="5:pRR1zhQ th7);RRh:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRVRHR=pRR0)RE
CMRRRRRCRs0MksR''4;R
RRDRC#RC
RRRRR0sCkRsM';j'
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?=;R

RR--QR8:BU3(
VRRk0MOHRFM""?=RR5p:QR1t7h ;RR):hRQa  t)s2RCs0kMQRAa#RH
LRRCMoH
RRRRRHVpRR=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;="
R
R-=-R=========================================================================
==
-RR-8RQ:3RB(Rg
RMVkOF0HM?R"/R="5Rp,)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR/=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?"/=;R

RR--QR8:Bj3U
VRRk0MOHRFM"=?/"pR5,RR):QR1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR/=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?"/=;R

RR--QR8:B43U
VRRk0MOHRFM"=?/"pR5Rh:Rq)azqRp;)RR:zQh1t7h 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR/=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?"/=;R

RR--QR8:B.3U
VRRk0MOHRFM"=?/"pR5RQ:Rhta  R);)RR:1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRVRHR/pR=RR)0MEC
RRRRsRRCs0kM4R''R;
RCRRD
#CRRRRRCRs0MksR''j;R
RRMRC8VRH;R
RCRM8VOkM0MHFR/"?=
";
-RR-8RQ:3RBURd
RMVkOF0HM?R"/R="5:pRR1zhQ th7);RRh:Rq)azqRp2skC0sAMRQHaR#R
RLHCoMR
RRVRHR/pR=RR)0MEC
RRRRsRRCs0kM4R''R;
RCRRD
#CRRRRRCRs0MksR''j;R
RRMRC8VRH;R
RCRM8VOkM0MHFR/"?=
";
-RR-8RQ:3RBURc
RMVkOF0HM?R"/R="5:pRRt1Qh; 7R:)RRaQh )t 2CRs0MksRaAQR
H#RCRLo
HMRRRRHpVRRR/=)ER0CRM
RRRRR0sCkRsM';4'
RRRR#CDCR
RRRRRskC0s'MRj
';RRRRCRM8H
V;RMRC8kRVMHO0F"MR?"/=;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1(34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413(R
RVOkM0MHFRD"#N5"RqR)t:hRz1hQt R7;BhmzaRR:Q hat2 )R0sCkRsMzQh1t7h R
H#RCRLo
HMRRRRH5VRBhmza=R>RRj20MEC
RRRRsRRCs0kM]R1Q_wapa w5tq),mRBz2ha;R
RRDRC#RC
RRRRR0sCkRsM1w]QaQ_)t5]aq,)tRm-Bz2ha;R
RRMRC8VRH;R
RCRM8VOkM0MHFRD"#N
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14HUR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4URkRVMHO0F"MR#"DNR)5qtRR:1hQt R7;BhmzaRR:Q hat2 )R0sCkRsM1hQt H7R#R
RLHCoMR
RRVRHRm5BzRha>j=R2ER0CRM
RRRRR0sCkRsM1w]Qa _pwqa5)Rt,Bhmza
2;RRRRCCD#
RRRRsRRCs0kM]R1Q_wa)]Qta)5qt-,RBhmza
2;RRRRCRM8H
V;RMRC8kRVMHO0F"MR#"DN;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1g34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413gR
RVOkM0MHFRs"#N5"RqR)t:hRz1hQt R7;BhmzaRR:Q hat2 )R0sCkRsMzQh1t7h R
H#RCRLo
HMRRRRH5VRBhmza=R>RRj20MEC
RRRRsRRCs0kM]R1Q_wa)]Qta)5qtB,Rmazh2R;
RCRRD
#CRRRRRCRs0MksRQ1]wpa_ 5waq,)tRm-Bz2ha;R
RRMRC8VRH;R
RCRM8VOkM0MHFRs"#N
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R1.HjR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
.jRkRVMHO0F"MR#"sNR)5qtRR:1hQt R7;BhmzaRR:Q hat2 )R0sCkRsM1hQt H7R#R
RLHCoMR
RRVRHRm5BzRha>j=R2ER0CRM
RRRRR0sCkRsM1w]QaQ_)t5]aq,)tRzBmh;a2
RRRR#CDCR
RRRRRskC0s1MR]aQw_wp a)5qt-,RBhmza
2;RRRRCRM8H
V;RMRC8kRVMHO0F"MR#"sN;R

RMVkOF0HMmRa_1zhQ th7qR5):tRRahqzp)q;QR1Z) _ :1RR1zhQ th7R2
RsRRCs0kMhRz1hQt H7R#R
RLHCoMR
RRCRs0MksR_amzQh1t7h R)5qt=RR>)RqtR,
RRRRRRRRRRRRRRRRRRRRR1RRQRZ =1>RQ_Z )' 1DoCM0;E2
CRRMV8Rk0MOHRFMazm_ht1Qh; 7
R
RVOkM0MHFR_am1hQt 57RqR)t:hRQa  t)1;RQ_Z )R 1:QR1t7h 2R
RRCRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMmRa_t1QhR 75tq)R>R=Rtq),R
RRRRRRRRRRRRRRRRRRRRR1 QZRR=>1 QZ_1) 'MDCo20E;R
RCRM8VOkM0MHFR_am1hQt 
7;
VRRk0MOHRFM)Q 1Z5 Rq,)tRZ1Q  _)1RR:zQh1t7h 2R
RRCRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsM)Q 1Z5 RqR)tRRRRRR=>q,)t
RRRRRRRRRRRRRRRRRRRh_ W1 QZRR=>1 QZ_1) 'MDCo20E;R
RCRM8VOkM0MHFR1) Q;Z 
R
RVOkM0MHFR1) QRZ 5tq),QR1Z) _ :1RRt1Qh2 7
RRRR0sCkRsM1hQt H7R#R
RLHCoMR
RRCRs0MksR1) QRZ 5tq)RRRRR>R=Rtq),R
RRRRRRRRRRRRRRRRRRWh _Z1Q >R=RZ1Q  _)1C'DMEo02R;
R8CMRMVkOF0HM R)1 QZ;R

RR--QR8:p634RR
RVOkM0MHFRM"N85"RpRR:A;QaR:)RR1zhQ th7s2RCs0kMhRz1hQt H7R#R
RLHCoMR
RRCRs0MksR1zhQ th7pR5R8NMRaAQ_Be a5m));22
CRRMV8Rk0MOHRFM"8NM"
;
R-R-R:Q8R4p3nRR
RMVkOF0HMNR"MR8"5:pRR1zhQ th7);RRA:RQRa2skC0szMRht1QhR 7HR#
RoLCHRM
RsRRCs0kMhRz1hQt 57RA_Qaea Bmp)52MRN82R);R
RCRM8VOkM0MHFRM"N8
";
-RR-8RQ:3Rp4
(RRkRVMHO0F"MRFRs"5:pRRaAQ;RR):hRz1hQt R72skC0szMRht1QhR 7HR#
RoLCHRM
RsRRCs0kMhRz1hQt 57RpsRFRaAQ_Be a5m));22
CRRMV8Rk0MOHRFM""Fs;R

RR--QR8:pU34RR
RVOkM0MHFRs"F"pR5Rz:Rht1Qh; 7R:)RRaAQ2CRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h RQ5Aa _eB)am5Rp2F)sR2R;
R8CMRMVkOF0HMFR"s
";
-RR-8RQ:3Rp4
gRRkRVMHO0F"MRM8NM"pR5RA:RQRa;)RR:zQh1t7h 2CRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h RR5pM8NMRaAQ_Be a5m));22
CRRMV8Rk0MOHRFM"MMN8
";
-RR-8RQ:3Rp.
jRRkRVMHO0F"MRM8NM"pR5Rz:Rht1Qh; 7R:)RRaAQ2CRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h RQ5Aa _eB)am5Rp2M8NMR;)2
CRRMV8Rk0MOHRFM"MMN8
";
-RR-8RQ:3Rp.
4RRkRVMHO0F"MRM"FsRR5p:QRAa);RRz:Rht1Qh2 7R0sCkRsMzQh1t7h R
H#RCRLo
HMRRRRskC0szMRht1QhR 75MpRFAsRQea_ mBa)25)2R;
R8CMRMVkOF0HMMR"F;s"
R
R-Q-R8p:R3R..
VRRk0MOHRFM"sMF"pR5Rz:Rht1Qh; 7R:)RRaAQ2CRs0MksR1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMzQh1t7h RQ5Aa _eB)am5Rp2MRFs)
2;RMRC8kRVMHO0F"MRM"Fs;R

RR--QR8:pd3.RR
RVOkM0MHFRF"Gs5"RpRR:A;QaR:)RR1zhQ th7s2RCs0kMhRz1hQt H7R#R
RLHCoMR
RRCRs0MksR1zhQ th7pR5RsGFRaAQ_Be a5m));22
CRRMV8Rk0MOHRFM"sGF"
;
R-R-R:Q8R.p3cRR
RMVkOF0HMGR"FRs"5:pRR1zhQ th7);RRA:RQRa2skC0szMRht1QhR 7HR#
RoLCHRM
RsRRCs0kMhRz1hQt 57RA_Qaea Bmp)52FRGs2R);R
RCRM8VOkM0MHFRF"Gs
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3Rp.H6R#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3R.6
VRRk0MOHRFM"FGMs5"RpRR:A;QaR:)RR1zhQ th7s2RCs0kMhRz1hQt H7R#R
RLHCoMR
RRCRs0MksR1zhQ th7pR5RFGMsQRAa _eB)am52)2;R
RCRM8VOkM0MHFRM"GF;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3R.nHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:pn3.RR
RVOkM0MHFRM"GFRs"5:pRR1zhQ th7);RRA:RQRa2skC0szMRht1QhR 7HR#
RoLCHRM
RsRRCs0kMhRz1hQt 57RA_Qaea Bmp)52MRGF)sR2R;
R8CMRMVkOF0HMGR"M"Fs;R

RR--QR8:p(3.RR
RVOkM0MHFRM"N85"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt H7R#R
RLHCoMR
RRCRs0MksRt1QhR 75NpRMA8RQea_ mBa)25)2R;
R8CMRMVkOF0HMNR"M;8"
R
R-Q-R8p:R3R.U
VRRk0MOHRFM"8NM"pR5R1:RQ th7);RRA:RQRa2skC0s1MRQ th7#RH
LRRCMoH
RRRR0sCkRsM1hQt 57RA_Qaea Bmp)52MRN82R);R
RCRM8VOkM0MHFRM"N8
";
-RR-8RQ:3Rp.
gRRkRVMHO0F"MRFRs"5:pRRaAQ;RR):QR1t7h 2CRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMQR1t7h RR5pFAsRQea_ mBa)25)2R;
R8CMRMVkOF0HMFR"s
";
-RR-8RQ:3Rpd
jRRkRVMHO0F"MRFRs"5:pRRt1Qh; 7R:)RRaAQ2CRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMQR1t7h RQ5Aa _eB)am5Rp2F)sR2R;
R8CMRMVkOF0HMFR"s
";
-RR-8RQ:3Rpd
4RRkRVMHO0F"MRM8NM"pR5RA:RQRa;)RR:1hQt R72skC0s1MRQ th7#RH
LRRCMoH
RRRR0sCkRsM1hQt 57RpNRMMA8RQea_ mBa)25)2R;
R8CMRMVkOF0HMMR"N"M8;R

RR--QR8:p.3dRR
RVOkM0MHFRN"MMR8"5:pRRt1Qh; 7R:)RRaAQ2CRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMQR1t7h RQ5Aa _eB)am5Rp2M8NMR;)2
CRRMV8Rk0MOHRFM"MMN8
";
-RR-8RQ:3Rpd
dRRkRVMHO0F"MRM"FsRR5p:QRAa);RR1:RQ th7s2RCs0kMQR1t7h R
H#RCRLo
HMRRRRskC0s1MRQ th7pR5RsMFRaAQ_Be a5m));22
CRRMV8Rk0MOHRFM"sMF"
;
R-R-R:Q8Rdp3cRR
RMVkOF0HMMR"FRs"5:pRRt1Qh; 7R:)RRaAQ2CRs0MksRt1QhR 7HR#
RoLCHRM
RsRRCs0kMQR1t7h RQ5Aa _eB)am5Rp2MRFs)
2;RMRC8kRVMHO0F"MRM"Fs;R

RR--QR8:p63dRR
RVOkM0MHFRF"Gs5"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt H7R#R
RLHCoMR
RRCRs0MksRt1QhR 75GpRFAsRQea_ mBa)25)2R;
R8CMRMVkOF0HMGR"F;s"
R
R-Q-R8p:R3Rdn
VRRk0MOHRFM"sGF"pR5R1:RQ th7);RRA:RQRa2skC0s1MRQ th7#RH
LRRCMoH
RRRR0sCkRsM1hQt 57RA_Qaea Bmp)52FRGs2R);R
RCRM8VOkM0MHFRF"Gs
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpdH(R#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3Rd(
VRRk0MOHRFM"FGMs5"RpRR:A;QaR:)RRt1Qh2 7R0sCkRsM1hQt H7R#R
RLHCoMR
RRCRs0MksRt1QhR 75GpRMRFsA_Qaea Bm))52
2;RMRC8kRVMHO0F"MRGsMF"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRdp3U#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3Rpd
URRkRVMHO0F"MRGsMF"pR5R1:RQ th7);RRA:RQRa2skC0s1MRQ th7#RH
LRRCMoH
RRRR0sCkRsM1hQt 57RA_Qaea Bmp)52MRGF)sR2R;
R8CMRMVkOF0HMGR"M"Fs;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpg3dRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rdp3gR
RVOkM0MHFRM"N85"RpRR:1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksR8NMRQ5Aa _eB)amR25p2R;
R8CMRMVkOF0HMNR"M;8"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RcjHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pj3c
VRRk0MOHRFM"8NM"pR5Rz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMMRN8AR5Qea_ mBa)pR52
2;RMRC8kRVMHO0F"MRN"M8;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp43cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp34R
RVOkM0MHFRN"MMR8"5:pRRt1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMNRMM58RA_Qaea Bm5)Rp;22
CRRMV8Rk0MOHRFM"MMN8
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcH.R#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
c.RkRVMHO0F"MRM8NM"pR5Rz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMNRMM58RA_Qaea Bm5)Rp;22
CRRMV8Rk0MOHRFM"MMN8
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHdR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cdRkRVMHO0F"MRFRs"5:pRRt1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMsRFRQ5Aa _eB)amR25p2R;
R8CMRMVkOF0HMFR"s
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHcR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
ccRkRVMHO0F"MRFRs"5:pRR1zhQ th7s2RCs0kMQRAa#RH
LRRCMoH
RRRR0sCkRsMF5sRA_Qaea Bm5)Rp;22
CRRMV8Rk0MOHRFM""Fs;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp63cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp36R
RVOkM0MHFRF"Ms5"RpRR:1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksRsMFRQ5Aa _eB)amR25p2R;
R8CMRMVkOF0HMMR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RcnHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pn3c
VRRk0MOHRFM"sMF"pR5Rz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMFRMsAR5Qea_ mBa)pR52
2;RMRC8kRVMHO0F"MRM"Fs;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp(3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3(R
RVOkM0MHFRF"Gs5"RpRR:1hQt R72skC0sAMRQHaR#R
RLHCoMR
RRCRs0MksRsGFRQ5Aa _eB)amR25p2R;
R8CMRMVkOF0HMGR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RcUHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pU3c
VRRk0MOHRFM"sGF"pR5Rz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMFRGsAR5Qea_ mBa)pR52
2;RMRC8kRVMHO0F"MRG"Fs;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpg3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3gR
RVOkM0MHFRM"GFRs"5:pRRt1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMMRGF5sRA_Qaea Bm5)Rp;22
CRRMV8Rk0MOHRFM"FGMs
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3Rp6HjR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
6jRkRVMHO0F"MRGsMF"pR5Rz:Rht1Qh2 7R0sCkRsMARQaHR#
RoLCHRM
RsRRCs0kMMRGF5sRA_Qaea Bm5)Rp;22
CRRMV8Rk0MOHRFM"FGMs
";
-RR-=R==========================================================================R=
RR--#H0sMOoRFCMPsF#HMMRN8sRIHR0CFsbCNF0HMR#
RR--============================================================================

RRRkRVMHO0F0MRF0_#soHMRN5PDRkCRRRR:MRHR1zhQ th7s2RCs0kMaR1)tQhR
H#RRRRNNDH#PRHNCDkRRRR:hRz1hQt 475RR0FPkNDCC'DMEo02#RHRDPNk
C;RRRRPHNsNCLDR#sCkRD0:aR1)tQh504RFNRPD'kCDoCM0;E2
FSOMN#0Mh0RzR1R:aR1)tQh50.RF2R4RR:=5EF0CRs#='>RR;'2RRRRRR--MDkDRs#0H
MoSoLCHRM
RHRRVNRPD'kCDoCM0<ERR04RE
CMRRRRRCRs0MksR1hz;R
RRDRC#RC
RRRRRsVFRHHRMPRHNCDk'MsNoDCRF
FbSRRRRVRHRe5HNCDk5RH2=jR''02RE
CMSsSSCD#k025HRR:=';j'
RSSCCD#
RSSRsRRCD#k025HRR:=';4'
RSSCRM8H
V;RRRRRMRC8FRDF
b;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_0MsHoR;
RR
RVOkM0MHFR_0F#H0sM5oRPkNDCRRRRRR:H1MRQ th7s2RCs0kMaR1)tQhR
H#RRRRNNDH#PRHNCDkRRRR:QR1t7h 504RFNRPD'kCDoCM0RE2HP#RNCDk;R
RRNRPsLHNDsCRCD#k0RR:1Qa)h4t5RR0FPkNDCC'DMEo02S;
O#FM00NMR1hzRRR:1Qa)h.t5RR0F4:2R=FR50sEC#>R=R''R2R;RR-RR-kRMD#DR0MsHoR
RLHCoMR
RRVRHRDPNkDC'C0MoERR<4ER0CRM
RRRRR0sCkRsMh;z1
RRRR#CDCR
RRRRRVRFsHMRHRNHPD'kCsoNMCFRDFRb
RRRRRRRRH5VRHDeNkHC52RR='2j'RC0EMS
SS#sCk5D0H:2R=jR''S;
SDRC#SC
SRRRR#sCk5D0H:2R=4R''S;
SMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_s#0H;Mo

RRRkRVMHO0F0MRF#_F0MsHoPR5NCDkRz:Rht1Qh2 7R0sCkRsM1Qa)hHtR#R
RLHCoMR
RRCRs0MksR_0FFs#0H5MoA_Qaea Bm5)RPkNDC;22
CRRMV8Rk0MOHRFM0FF_#H0sM
o;
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:1hQt R72skC0s1MRah)Qt#RH
RRRRMOF#M0N0CRs#0kD_MDCoR0E:hRQa  t)=R:RN5PD'kCDoCM0.E+2;/d
RRRRMOF#M0N0NRb8RRRRRRRRRRR:QRAa _eB)am504RFsR5CD#k0C_DMEo0*-dRRDPNkDC'C0MoE
22RRRRR=R:R05FE#CsRR=>PkNDCPR5NCDk'VDC0;22R-R-R0 GCRM8#MHoR0LH
LRRCMoH
RRRR0sCkRsM0FF_#H0sMbo5N&8RRaAQ_Be aRm)5DPNk2C2;R
RCRM8VOkM0MHFR_0FFs#0H;Mo
R
RVOkM0MHFR_0FEs#0HRMo5DPNk:CRR1zhQ th7s2RCs0kMaR1)tQhR
H#RCRLo
HMRRRRskC0s0MRF#_E0MsHoQ5Aa _eB)amRN5PD2kC2R;
R8CMRMVkOF0HMFR0_0E#soHM;R

RMVkOF0HMFR0_0E#soHMRN5PDRkC:QR1t7h 2CRs0MksR)1aQRhtHR#
RORRF0M#NRM0skC#DD0_C0MoERR:Q hatR ):5=RPkNDCC'DMEo0+/d2cR;
RORRF0M#NRM0bRN8RRRRRRRRRRR:A_Qaea Bm4)5RR0F5#sCk_D0DoCM0cE*RP-RNCDk'MDCo20E2R
RRRRR:5=RFC0Es=#R>NRPDRkC5DPNkDC'C2V02R;R- -RGM0C8HR#oLMRHR0
RoLCHRM
RsRRCs0kMFR0_0E#soHM58bNRA&RQea_ mBa)PR5NCDk2
2;RMRC8kRVMHO0F0MRF#_E0MsHoR;
RM
C8zRhvQ )BQ_Aa
;

