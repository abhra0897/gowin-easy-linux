`define getname(oriName,tmodule_name) \~oriName.tmodule_name 

`ifdef CONST_VH
`else
`define CONST_VH

`define	PRODUCT_ID			32'h00021009

`ifdef ADDR_WIDTH_24
`define	ADDR_MSB			23
`define SLV_OFFSET_UNIT		10
`else
`define	ADDR_MSB			31
`define SLV_OFFSET_UNIT		20
`endif

`define SPACE_MSB			(`ADDR_DECODE_WIDTH - 1)

`define SLV_0

`ifdef ADDR_WIDTH_24
`define SLV0_SIZE			3
`else
`define SLV0_SIZE			1
`endif

`ifndef SLV0_OFFSET
`define	SLV0_OFFSET		`ADDR_DECODE_WIDTH'h0
`endif

`define SLV0_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV0_SIZE - 1)
`define SLV1_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV1_SIZE - 1)
`define SLV2_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV2_SIZE - 1)
`define SLV3_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV3_SIZE - 1)
`define SLV4_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV4_SIZE - 1)
`define SLV5_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV5_SIZE - 1)
`define SLV6_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV6_SIZE - 1)
`define SLV7_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV7_SIZE - 1)
`define SLV8_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV8_SIZE - 1)
`define SLV9_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV9_SIZE - 1)
`define SLV10_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV10_SIZE - 1)
`define SLV11_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV11_SIZE - 1)
`define SLV12_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV12_SIZE - 1)
`define SLV13_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV13_SIZE - 1)
`define SLV14_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV14_SIZE - 1)
`define SLV15_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV15_SIZE - 1)
`define SLV16_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV16_SIZE - 1)
`define SLV17_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV17_SIZE - 1)
`define SLV18_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV18_SIZE - 1)
`define SLV19_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV19_SIZE - 1)
`define SLV20_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV20_SIZE - 1)
`define SLV21_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV21_SIZE - 1)
`define SLV22_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV22_SIZE - 1)
`define SLV23_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV23_SIZE - 1)
`define SLV24_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV24_SIZE - 1)
`define SLV25_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV25_SIZE - 1)
`define SLV26_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV26_SIZE - 1)
`define SLV27_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV27_SIZE - 1)
`define SLV28_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV28_SIZE - 1)
`define SLV29_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV29_SIZE - 1)
`define SLV30_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV30_SIZE - 1)
`define SLV31_OFFSET_LSB		(`SLV_OFFSET_UNIT + `SLV31_SIZE - 1)
`define OFFSET_MSB			`SPACE_MSB


`define SLV1_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV1_OFFSET} | 33'd`SLV1_SIZE)
`define SLV2_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV2_OFFSET} | 33'd`SLV2_SIZE)
`define SLV3_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV3_OFFSET} | 33'd`SLV3_SIZE)
`define SLV4_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV4_OFFSET} | 33'd`SLV4_SIZE)
`define SLV5_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV5_OFFSET} | 33'd`SLV5_SIZE)
`define SLV6_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV6_OFFSET} | 33'd`SLV6_SIZE)
`define SLV7_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV7_OFFSET} | 33'd`SLV7_SIZE)
`define SLV8_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV8_OFFSET} | 33'd`SLV8_SIZE)
`define SLV9_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV9_OFFSET} | 33'd`SLV9_SIZE)
`define SLV10_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV10_OFFSET} | 33'd`SLV10_SIZE)
`define SLV11_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV11_OFFSET} | 33'd`SLV11_SIZE)
`define SLV12_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV12_OFFSET} | 33'd`SLV12_SIZE)
`define SLV13_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV13_OFFSET} | 33'd`SLV13_SIZE)
`define SLV14_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV14_OFFSET} | 33'd`SLV14_SIZE)
`define SLV15_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV15_OFFSET} | 33'd`SLV15_SIZE)
`define SLV16_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV16_OFFSET} | 33'd`SLV16_SIZE)
`define SLV17_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV17_OFFSET} | 33'd`SLV17_SIZE)
`define SLV18_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV18_OFFSET} | 33'd`SLV18_SIZE)
`define SLV19_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV19_OFFSET} | 33'd`SLV19_SIZE)
`define SLV20_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV20_OFFSET} | 33'd`SLV20_SIZE)
`define SLV21_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV21_OFFSET} | 33'd`SLV21_SIZE)
`define SLV22_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV22_OFFSET} | 33'd`SLV22_SIZE)
`define SLV23_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV23_OFFSET} | 33'd`SLV23_SIZE)
`define SLV24_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV24_OFFSET} | 33'd`SLV24_SIZE)
`define SLV25_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV25_OFFSET} | 33'd`SLV25_SIZE)
`define SLV26_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV26_OFFSET} | 33'd`SLV26_SIZE)
`define SLV27_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV27_OFFSET} | 33'd`SLV27_SIZE)
`define SLV28_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV28_OFFSET} | 33'd`SLV28_SIZE)
`define SLV29_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV29_OFFSET} | 33'd`SLV29_SIZE)
`define SLV30_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV30_OFFSET} | 33'd`SLV30_SIZE)
`define SLV31_CFG_REG		({{33-`ADDR_DECODE_WIDTH{1'b0}}, `SLV31_OFFSET} | 33'd`SLV31_SIZE)
`define REG_ADDR_WIDTH		8
`define	REG_ADDR_MSB		(`REG_ADDR_WIDTH + 1)

`endif
