--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..4N/OGlbNbC/s#GHHDMDG/HoL/C#M_b0NsN/MdsMNl_Is_38PEyf4R

--

-----
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFR0LFECRsNN8RMI8RsCH0
R--aoNsC:0RRDXHH
MG---
-jR4/Rj41RC0Wa)Q m_v7q _Rs5IHR0Cb0Fs2FR0Rq) 7Q_w)R1aH8MRCkVNDV0RF-s
-RRROVFMD0HOR#sCF0DkHRFMbbksF3#CRV)CC0sRFHResG0C-RQQwqutRM]N8FLF	-
-RBRRE0NbCRs."Hz#MAoRD	FORD1CC)O0qvvRCslF$#"RCHO0F
M3
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)v)h__HWR#o
SCsMCH5OR
RSRRNRVl$HDR#:R0MsHo=R:RF"MM;C"
ISSHE80RH:RMo0CC:sR=;R4RS
SNs88I0H8ERR:HCM0oRCs:n=R;RRRRRRRRR--LRHoCkMFoVERF8sRCEb0
8SSCEb0RH:RMo0CC:sR=URc;S
S80Fk_osCRL:RFCFDN:MR=NRVD;#CRRRRR-R-R#ENR0FkbRk0s
CoSHS8MC_soRR:LDFFCRNM:V=RNCD#;RRRRRRRRR--ERN#8NN0RbHMks0RCRo
RRRRRsRR#80_NR0N:0R#soHM;S
SIls_F:8CRs#0HRMo:"=RWa)Q Q_w)"1a;S
Ss8N8sC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#CRsNN8R8C8s#s#RCSo
S8IN8ss_C:oRRFLFDMCNR=R:RDVN#RCRRRRR-E-RNI#RsCH0R8N8s#C#RosC
2SS;b
SFRs05S
S7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
S)7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2S;
Sh7QRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7Wq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;S SWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlSpSBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMSBSmp:iRRRHM#_08DHFoOR;RRRRR-F-RbO0RD	FORsVFR8I_F
k0RRRRRRRR :hRRRHM#_08DHFoOR;RRRRRR-R-RNCML
DCRRRRRRRRWh_ RH:RM0R#8F_Do;HORRRRRRRR-C-RMDNLCR
RRRRRR1R)aRR:H#MR0D8_FOoHRRRRRRRR-#-R#Rs
RRRRR2RR;M
C8MRC0$H0Rv)qh__)W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCLODF	N_slVRFRv)qh__)W#RH
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks5F"hRNsC8s/IHR0COVFMD0HORCOEOR	31kHlDHN0FlMRHN#l0ROEb#F#HCLDR"!!2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
CRRMo8RCC0_M88_CEb0;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHo-;
-0N0skHL0oCRCsMCNs0F_bsCFRs0FLVRD	FO_lsNRN:RsHOE00COkRsCHV#Rk_MOH0MH58sN8ss_C;o2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFM#H0sM#o.DNP5R#:R0MsHos2RCs0kM0R#8F_Do_HOP0COFHsR#N
PsLHND#CRD:PRR8#0_oDFHPO_CFO0s'5NEEHo-DN'F8IRF0IMF2Rj;N
PsLHNDHCRRH:RMo0CC
s;LHCoMR
RVRFsHMRHR0jRFDR#PH'EoDERF
FbRRRRH5VRN'5NEEHo-RH2=4R''02RE
CMS#RRDHP52=R:R''4;C
SD
#CS#RRDHP52=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#;DP
8CMRs#0H.Mo#;DP
MVkOF0HMDR#P0.#soHM5:NRR8#0_oDFHPO_CFO0ss2RCs0kM0R#soHMR
H#PHNsNCLDR:#RRs#0H5MoNH'EoNE-'IDF+84RF0IMF2R4;N
PsLHNDHCRRH:RMo0CC
s;LHCoMR
RVRFsHMRHRDN'F0IRF'RNEEHoRFDFbR
RRVRHR55NH=2RR''42ER0CSM
R5R#H'-ND+FI4:2R=4R''S;
CCD#
RSR#-5HNF'DI2+4RR:=';j'
MSC8VRH;R
RCRM8DbFF;R
RskC0s#MR;M
C8DR#P0.#soHM;0
N0LsHkR0CGbO_s#FbR#:R0MsHo-;
-MOF#M0N0sR#PRND:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2RjRR:=#H0sM#o.DsP5#80_N20N;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFR0oC_FOEH_OCI0H8EH5I8R0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;N
PsLHND8CRH.Pd,HR8P,4nRP8HU8,RH,PcRP8H.8,RHRP4:MRH0CCosL;
CMoH
8RRH.PdRR:=58IH04E-2n/d;R
R84HPn=R:RH5I8-0E442/UR;
RP8HU=R:RH5I8-0E4g2/;R
R8cHPRR:=58IH04E-2;/c
8RRHRP.:5=RI0H8E2-4/
.;RHR8P:4R=IR5HE80-;42
HRRV8R5HRP4>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>.RRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HcRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8UHPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HnP4Rj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
R--RRHV5P8Hd>.RRRj20MEC
R--RPRRN:DR=NRPDRR+4-;
-CRRMH8RVR;
RRHV5DPNR.>R2ER0CRM
RsRRCs0kM.R5RR**PRND+RR.*5*RPRND-2Rd2R;
R#CDCR
RRCRs0MksRR5.*P*RN;D2
CRRMH8RVC;
Mo8RCO0_EOFHCH_I8;0E
MVkOF0HMCRo0E_OFCHO_b8C08E5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHND8CR_FOEH_OC80CbERR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E>4RUgR.20MEC
RRRRO8_EOFHCC_8bR0E:4=RncdU;R
RCHD#V8R5CEb0RR<=U.4gR8NMRb8C0>ERRgcjnRR20MEC
RRRRO8_EOFHCC_8bR0E:U=R4;g.
CRRDV#HRC58bR0E<c=RjRgnNRM880CbERR>.Ujc2ER0CRM
R8RR_FOEH_OC80CbE=R:RgcjnR;
R#CDH5VR80CbE=R<Rc.jUMRN8CR8bR0E>jR4.2cRRC0EMR
RR_R8OHEFO8C_CEb0RR:=.Ujc;R
RCHD#V8R5CEb0RR<=4cj.R8NMRb8C0>ERR.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.4jcR;
R#CDH5VR80CbE=R<R.642ER0CRM
R8RR_FOEH_OC80CbE=R:R.64;R
RCRM8H
V;RCRs0MksRO8_EOFHCC_8b;0E
8CMR0oC_FOEH_OC80CbEV;
k0MOHRFMo_C0I0H8EF_l85_UOHEFOIC_8RR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCI0H8EF_l8R_U:MRH0CCosL;
CMoH
HRRVOR5EOFHC8_IRU>R2ER0CRM
RIRRHE80_8lF_:UR=EROFCHO_RI8-OR5EOFHC8_IR8lFR;U2
CRRD
#CRRRRI0H8EF_l8R_U:O=REOFHC8_I;R
RCRM8H
V;RCRs0MksR8IH0lE_FU8_;M
C8CRo0H_I8_0El_F8U
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R0oC_FOEH_OCI0H8EH5I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:4=RncdU/0oC_8IH0lE_FU8_5OI_EOFHCH_I820E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:o=RCO0_EOFHCC_8b50E80CbE
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:Rn54d/Uc8E_OFCHO_b8C0RE2+5R54Undc_/8OHEFO8C_CEb02RR/U
2;
MVkOF0HMCRo0k_MlC_OD5D#I:8RR0HMCsoC;FOEH_OCI:8RR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRlMk_DOCD:#RR0HMCsoC;C
Lo
HMRkRMlC_ODRD#:5=RI48-2E/OFCHO_RI8+;R4
sRRCs0kMkRMlC_OD;D#
8CMR0oC_lMk_DOCD
#;
MVkOF0HMCRo0H_#xIC5M:ORR0HMCsoC;MR8ORR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
RRRskC0sIMRM*ORRO8M;M
C8CRo0H_#x
C;
MVkOF0HMCRo0F_LF5D88H_#x:CRR0HMCsoC;_RI#CHxRH:RMo0CCRs;8I_ORH:RMo0CCRs;II_ORH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMH5VR8H_#x<CR=_RI#CHx2ER0CRM
R0sCkRsM8I_O;D
C#RC
R0sCkRsMII_O;M
C8VRH;M
C8CRo0F_LF;D8
F
OMN#0MO0REOFHCH_I8R0E:MRH0CCos=R:R0oC_FLFDo85C#0_H5xCo_C0M_klODCD#H5I8,0ERO8_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_R8OHEFO8C_CEb02
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSS_R8OHEFOIC_HE80,_RIOHEFOIC_HE802O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:R0oC_FLFDo85C#0_H5xCo_C0M_klODCD#H5I8,0ERO8_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_R8OHEFO8C_CEb02
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRo_C0#CHx50oC_lMk_DOCDI#5HE80,_RIOHEFOIC_HE802C,o0k_MlC_OD5D#80CbEI,R_FOEH_OC80CbE,22
SSSSSSSSSSSRRRR58IH04E-2_/8OHEFOIC_HE80,IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSR5RR80CbE2-4/O8_EOFHCC_8b,0ERC58b-0E4I2/_FOEH_OC80CbE+2RRS4;RF
OMN#0Mx0RCRsF:0R#8F_Do_HOP0COFOs5EOFHCH_I8*0EI0H8Ek_MlC_OD-D#I0H8ER-48MFI0jFR2=R:R05FE#CsRR=>'2j';F
OMN#0M#0RsDPN_P#DR#:R0D8_FOoH_OPC05FsOHEFOIC_HE80*8IH0ME_kOl_C#DD-84RF0IMF2RjRR:=xFCsR#&R0MsHoD.#P#5s0N_80;N2
MOF#M0N0sR#PRND:0R#soHM5FOEH_OCI0H8EH*I8_0EM_klODCD#FR8IFM0RR42:#=RD#P.0MsHos5#P_ND#2DP;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L.k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#.:kRF0k_L#0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RUI0H8Ek_MlC_OD+D#(FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkURR:F_k0LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjd,R.H*I8_0EM_klODCD#4+dRI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Ldk#.RR:F_k0Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDkRF0C_so:4RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FOFEF#LCRCC0IC7MRQNhRMF8Rkk0b0VRFRFADO)	Rq#v
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqR)7
7)#MHoNIDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--s8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDqR)7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC)7q7)H
#oDMNR7Wq70)_l:bRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCRq)77
o#HMRND7_Qh0Rlb:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCQR7hH
#oDMNR_W 0Rlb:0R#8F_Do;HORRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDMWCR -
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0k_Mlc_n5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/;nc
HRRV5R580CbEFRl8cRn2RR>cRU20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FCds_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8cRn2C;
Mo8RCD0_CFV0P_Csd
.;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_nO;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5nc80CbE
2;O#FM00NMRVDC0CFPs._dRH:RMo0CC:sR=CRo0C_DVP0FCds_.C58b20E;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bCnRc#HN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._d##RHRsNsN5$RM_klODCD_Rd.8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bC4Rn#HN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#_c:#RR0Fk_#Lk_b0$Cc_n#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kd#_.:#RR0Fk_#Lk_b0$C._d#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_k4#_n:#RR0Fk_#Lk_b0$Cn_4#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNFDRkC0_M._dR#:R0D8_FOoH;H
#oDMNR0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDNRs8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDI_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDIN_s8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjjjjjjRj"&NRs8C_so25j;R
SRDRRFII_Ns88RR<="jjjjjjjjjjjjRj"&NRI8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjjjRj"&NRs8C_soR548MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjjRj"&NRI8C_soR548MFI0jFR2S;
CRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjjRj"&NRs8C_soR5.8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj&"RR8IN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjj"RR&s_N8s5CodFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=RjjjjjjjjjRj"&NRI8C_soR5d8MFI0jFR2S;
CRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80R6=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj"jjRs&RNs8_Cco5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjj"RR&I_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjj"RR&s_N8s5Co6FR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjjj&"RR8IN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjj"RR&s_N8s5ConFR8IFM0R;j2
DSSFII_Ns88RR<="jjjjjjj"RR&I_N8s5ConFR8IFM0R;j2
MSC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjjjjjRj"&NRs8C_soR5(8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjjj&"RR8IN_osC58(RF0IMF2Rj;C
SMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjRj"&NRs8C_soR5U8MFI0jFR2S;
SIDF_8IN8<sR=jR"jjjj"RR&I_N8s5CoUFR8IFM0R;j2
MSC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj&"RR8sN_osC58gRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjRj"&NRI8C_soR5g8MFI0jFR2S;
CRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RSRRFRDIN_s8R8s<"=Rj"jjRs&RNs8_C4o5jFR8IFM0R;j2
DSSFII_Ns88RR<="jjj"RR&I_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDIN_s8R8s<"=RjRj"&NRs8C_so454RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjRj"&NRI8C_so454RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R''jRs&RNs8_C4o5.FR8IFM0R;j2
DSSFII_Ns88RR<='Rj'&NRI8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FIs8N8s=R<R8sN_osC5R4d8MFI0jFR2S;
RRRRD_FII8N8s=R<R8IN_osC5R4d8MFI0jFR2S;
CRM8oCCMsCN0Rdz4;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR4Rzc:RRRRHV5M8H_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piRh7Q2CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2S;
CRM8oCCMsCN0R6z4;R

R7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRR4RnsRH:RVsR5Ns88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
R--RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
R--RRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMRFbsO#C#;-
-S8CMRMoCC0sNC4Rzn
s;-R-RR4Rz(:sRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)S;
CRM8oCCMsCN0Rnz4s
;
SR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoWB_mpRi
RzRR4RnIRH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4;nI
RRRR(z4IRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;C
SMo8RCsMCNR0CzI4(;R

R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141S4
zR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
RRRR4SzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24cRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.Rz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_ncdUXR47:NRDLRCDH"#RWa)Q m_v7q _=q) 7Q_w),1aRe1)qAp_=&"RRP#sN[D5+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUXR47:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4Undc&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424Undc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2S;
SCSLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4:7RRv)qA_4n114_4R
SRRRRRRRRRbRRFRs0lRNb5q7Q5Rj2=H>RMC_so25[,7Rq7R)q=D>RFII_Ns885R4d8MFI0jFR27,RQ=AR>jR""q,R7A7)RR=>D_FIs8N8sd54RI8FMR0Fj
2,SSSS Rhq=W>R_, hR)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=> Rh,1A1)RR=>),1aRAW RR=>',j'RiBpA>R=RpmBiS,
SRSRRmR7q>R=RCFbM7,RmjA52>R=R0Fk_#Lk4,5H[;22
R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRSRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1.1S.
zR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qvU.4gXR.7:NRDLRCDH"#RWa)Q m_v7q _=q) 7Q_w),1aRe1)qAp_=&"RRP#sN.D5*.[+RI8FMR0F.+*[4&2RRR",Wa)Q m_v7A _=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..X7RR:DCNLD#RHR7"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*UgR.2&WR""RR&HCM0o'CsHolNC*5[.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4U2*4,g.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;.2
SSSLHCoMR
RRRRRRRRRRARS)_qvU.4gXR.7:qR)vnA4__1.1S.
RRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7q7)RR=>D_FII8N8s.54RI8FMR0FjR2,7RQA=">Rj,j"R7q7)=AR>FRDIN_s858s48.RF0IMF2Rj,S
SSRRRRq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmp
i,SRSSR7RRm=qR>bRFCRM,75mA4=2R>kRF0k_L#H.5,[.*+,42RA7m5Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0RC
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R.2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzd;-
S-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:4RRRHV58N8s8IH0<ER=.R42CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;d4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gcjn7XcRD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5NDc+*[cFR8IFM0R[c*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgnc:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5cH*j2gnR"&RW&"RR0HMCsoC'NHlo[C5*Rc2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42cnjg,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*c;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
SSSSq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmp
i,SSSS7Rmq=F>Rb,CMRA7m5Rd2=F>RkL0_k5#cHc,R*d[+27,Rm.A52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSSA7m5R42=F>RkL0_k5#cH*,c[2+4,mR7A25jRR=>F_k0Lck#5RH,c2*[2R;
RRRRRRRRRRRRRFRRks0_Cco5*R[2<F=RkL0_k5#cH*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[4<2R=kRF0k_L#Hc5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R.2<F=RkL0_k5#cH*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+dRR<=F_k0Lck#5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1g1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv.UjcXRU7:NRDLRCDH"#RWa)Q m_v7q _=q) 7Q_w),1aRe1)qAp_=&"RRP#sNgD5*g[+RI8FMR0Fg+*[4&2RRR",Wa)Q m_v7A _=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUX7RR:DCNLD#RHR7"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*.cRU2&WR""RR&HCM0o'CsHolNC*5[g&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4.2*j,cURb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;g2
SSSLHCoMR
RRRRRRRRRRARS)_qv.UjcXRU7:qR)vnA4__1g1Rg
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77q>R=RIDF_8IN84s5jFR8IFM0R,j2RA7QRR=>"jjjjjjjjR",q)77A>R=RIDF_8sN84s5jFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25(RR=>F_k0LUk#5UH,*([+27,RmnA52>R=R0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R62=F>RkL0_k5#UH*,U[2+6,mR7A25cRR=>F_k0LUk#5UH,*c[+27,RmdA52>R=R0Fk_#LkU,5HU+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R.2=F>RkL0_k5#UH*,U[2+.,mR7A254RR=>F_k0LUk#5UH,*4[+27,RmjA52>R=R0Fk_#LkU,5HU2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ5uqj=2R>MRH_osC5[g*+,U2Ru7QA>R=R""j,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u=qR>bRFCRM,7Amu5Rj2=b>RN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d(
RRRRCRSMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_41U_4SU
zRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCR
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;cj
-S-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRcSz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;c4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_.4jcnX47RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5*4U[U+4RI8FMR0F4[U*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4Rn7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5H4cj.2RR&"RW"&MRH0CCosl'HN5oC[U*42RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*4.Rc,80CbER22&XR""RR&HCM0o'CsHolNC[55+*424;U2
SSSLHCoMR
RRRRRRRRRRARS)_qv4cj.X74nR):Rq4vAn4_1U4_1UR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7R)q=D>RFII_Ns8858gRF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sgFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A6542>R=R0Fk_#Lk4Hn5,*4n[6+427,Rm4A5c=2R>kRF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524dRR=>F_k0L4k#n,5H4[n*+24d,mR7A.542>R=R0Fk_#Lk4Hn5,*4n[.+427,Rm4A54=2R>kRF0k_L#54nHn,4*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524jRR=>F_k0L4k#n,5H4[n*+24j,mR7A25gRR=>F_k0L4k#n,5H4[n*+,g2RA7m5RU2=F>RkL0_kn#454H,n+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R(2=F>RkL0_kn#454H,n+*[(R2,75mAn=2R>kRF0k_L#54nHn,4*n[+27,Rm6A52>R=R0Fk_#Lk4Hn5,*4n[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmcA52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR7A25dRR=>F_k0L4k#n,5H4[n*+,d2RA7m5R.2=F>RkL0_kn#454H,n+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R42=F>RkL0_kn#454H,n+*[4R2,75mAj=2R>kRF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,QR7u=AR>jR"jR",7qmuRR=>FMbC,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RsbNH_0$L4k#n,5H.+*[4R2,7Amu5Rj2=b>RN0sH$k_L#54nH*,.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
RRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SSjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SSSSF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc;jN
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SS4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0CzNc4;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSScR.N:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_.64X7d.RD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5NDd[n*+Rdn8MFI0dFRn+*[4&2RRR",Wa)Q m_v7A _=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..Xd7RR:DCNLD#RHR7"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*6.&2RR""WRH&RMo0CCHs'lCNo5d[*n&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+462*4R.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42d;n2
SSSLHCoMR
RRRRRRRRRRRRRRRRRRRRRRRRRAv)q_.64X7d.R):Rq4vAnd_1nd_1nR
RRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmp
i,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,RmdA54=2R>kRF0k_L#5d.H.,d*d[+4R2,75mAdRj2=F>RkL0_k.#d5dH,.+*[d,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5g=2R>kRF0k_L#5d.H.,d*.[+gR2,75mA.RU2=F>RkL0_k.#d5dH,.+*[.,U2RA7m52.(RR=>F_k0Ldk#.,5Hd[.*+2.(,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rn2=F>RkL0_k.#d5dH,.+*[.,n2RA7m52.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR7Ac5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR7A.5.2>R=R0Fk_#LkdH.5,*d.[.+.27,Rm.A54=2R>kRF0k_L#5d.H.,d*.[+4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Aj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rm4A5g=2R>kRF0k_L#5d.H.,d*4[+gR2,75mA4RU2=F>RkL0_k.#d5dH,.+*[4,U2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5(=2R>kRF0k_L#5d.H.,d*4[+(R2,75mA4Rn2=F>RkL0_k.#d5dH,.+*[4,n2RA7m5246RR=>F_k0Ldk#.,5Hd[.*+246,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rc2=F>RkL0_k.#d5dH,.+*[4,c2RA7m524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7A.542>R=R0Fk_#LkdH.5,*d.[.+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5244RR=>F_k0Ldk#.,5Hd[.*+244,mR7Aj542>R=R0Fk_#LkdH.5,*d.[j+427,RmgA52>R=R0Fk_#LkdH.5,*d.[2+g,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAU=2R>kRF0k_L#5d.H.,d*U[+27,Rm(A52>R=R0Fk_#LkdH.5,*d.[2+(,mR7A25nRR=>F_k0Ldk#.,5Hd[.*+,n2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm6A52>R=R0Fk_#LkdH.5,*d.[2+6,mR7A25cRR=>F_k0Ldk#.,5Hd[.*+,c2RA7m5Rd2=F>RkL0_k.#d5dH,.+*[d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>F_k0Ldk#.,5Hd[.*+,.2RA7m5R42=F>RkL0_k.#d5dH,.+*[4R2,75mAj=2R>kRF0k_L#5d.H.,d*,[2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"7,RmRuq=F>Rb,CM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uAd=2R>NRbs$H0_#LkdH.5,[c*+,d2Ru7mA25.RR=>bHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>bHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>NRbs$H0_#LkdH.5,[c*2
2;RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S

SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;C

MN8RsHOE00COkRsCLODF	N_sl
;
NEsOHO0C0CksR_MFsOI_E	CORRFV)hqv_W)_R
H#VOkM0MHFRMVkOM_HHL05RL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
RRHV5RL20MEC
RRRR0sCk5sM"RhFs8CN/HIs0OCRFDMVHRO0OOEC	13RHDlkNF0HMHRl#0lNObERFH##LRDC!2!";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;RMRC8CRo0M_C8C_8b;0E
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;-
-Ns00H0LkCCRoMNCs0_FssFCbsF0RVFRM__sIOOEC	RR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFRs#0H.Mo#5DPNRR:#H0sMRo2skC0s#MR0D8_FOoH_OPC0RFsHP#
NNsHLRDC#RDP:0R#8F_Do_HOP0COFNs5'oEHE'-NDRFI8MFI0jFR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRMRRj0#FRDEP'HRoEDbFF
RRRRRHV5NN5'oEHE2-HR'=R4R'20MEC
RSR#5DPH:2R=4R''S;
CCD#
RSR#5DPH:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksRP#D;M
C80R#soHM.P#D;k
VMHO0F#MRD#P.0MsHoR5N:0R#8F_Do_HOP0COFRs2skC0s#MR0MsHo#RH
sPNHDNLCRR#:0R#soHM5EN'H-oENF'DIR+48MFI04FR2P;
NNsHLRDCHRR:HCM0o;Cs
oLCHRM
RsVFRHHRM'RNDRFI0NFR'oEHEFRDFRb
RHRRVNR55RH2=4R''02RE
CMS#RR5NH-'IDF+R42:'=R4
';S#CDCR
SRH#5-DN'F4I+2=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#C;
M#8RD#P.0MsHoN;
0H0sLCk0R_GObbsF#RR:#H0sM
o;-F-OMN#0M#0RsDPNR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2=R:Rs#0H.Mo#5DPs_#08NN02-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0E_OFCHO_8IH0IE5HE80RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jP;
NNsHLRDC8dHP.8,RHnP4,HR8PRU,8cHP,HR8PR.,84HPRH:RMo0CC
s;LHCoMR
R8dHP.=R:RH5I8-0E4d2/nR;
RP8H4:nR=IR5HE80-/424
U;RHR8P:UR=IR5HE80-/42gR;
RP8Hc=R:RH5I8-0E4c2/;R
R8.HPRR:=58IH04E-2;/.
8RRHRP4:5=RI0H8E2-4;R
RH5VR84HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRP.>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>cRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HURR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR84HPnRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;-
-RVRHRH58PRd.>2RjRC0EM-
-RRRRPRND:P=RN+DRR
4;-R-RCRM8H
V;RVRHRN5PDRR>.02RE
CMRRRRskC0s5MR.*R*RDPNR.+RRR**5DPNRd-R2
2;RDRC#RC
RsRRCs0kM.R5RR**P2ND;R
RCRM8H
V;CRM8o_C0OHEFOIC_HE80;k
VMHO0FoMRCO0_EOFHCC_8b50E80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDC8E_OFCHO_b8C0:ERR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RU>R42g.RC0EMR
RR_R8OHEFO8C_CEb0RR:=4UndcR;
R#CDH5VR80CbE=R<RgU4.MRN8CR8bR0E>jRcg2nRRC0EMR
RR_R8OHEFO8C_CEb0RR:=U.4g;R
RCHD#V8R5CEb0RR<=cnjgR8NMRb8C0>ERRc.jU02RE
CMRRRR8E_OFCHO_b8C0:ER=jRcg
n;RDRC#RHV5b8C0<ER=jR.cNURM88RCEb0R4>RjR.c2ER0CRM
R8RR_FOEH_OC80CbE=R:Rc.jUR;
R#CDH5VR80CbE=R<R.4jcMRN8CR8bR0E>4R6.02RE
CMRRRR8E_OFCHO_b8C0:ER=jR4.
c;RDRC#RHV5b8C0<ER=4R6.02RE
CMRRRR8E_OFCHO_b8C0:ER=4R6.R;
R8CMR;HV
sRRCs0kM_R8OHEFO8C_CEb0;M
C8CRo0E_OFCHO_b8C0
E;VOkM0MHFR0oC_8IH0lE_FU8_5FOEH_OCI:8RR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDR8IH0lE_FU8_RH:RMo0CC
s;LHCoMR
RH5VROHEFOIC_8RR>U02RE
CMRRRRI0H8EF_l8R_U:O=REOFHC8_IR5-ROHEFOIC_8FRl82RU;R
RCCD#
RRRR8IH0lE_FU8_RR:=OHEFOIC_8R;
R8CMR;HV
sRRCs0kMHRI8_0El_F8UC;
Mo8RCI0_HE80_8lF_
U;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=CRo0E_OFCHO_8IH0IE5HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=4UndcC/o0H_I8_0El_F8U_5IOHEFOIC_HE802O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=o_C0OHEFO8C_CEb05b8C0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=4R5ncdU/O8_EOFHCC_8b20ER5+R5d4nU8c/_FOEH_OC80CbE/2RR;U2
k
VMHO0FoMRCM0_kOl_C#DD5RI8:MRH0CCosE;OFCHO_RI8:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCkRMlC_ODRD#:MRH0CCosL;
CMoH
MRRkOl_C#DDRR:=5-I84O2/EOFHC8_IR4+R;R
RskC0sMMRkOl_C#DD;M
C8CRo0k_MlC_OD;D#
k
VMHO0FoMRC#0_H5xCIRMO:MRH0CCos8;RM:ORR0HMCsoC2CRs0MksR0HMCsoCR
H#LHCoMR
RR0sCkRsMIRMO*MR8OC;
Mo8RC#0_H;xC
k
VMHO0FoMRCL0_F8FD5#8_HRxC:MRH0CCosI;R_x#HCRR:HCM0o;CsRO8_IRR:HCM0o;CsROI_IRR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
RHV5#8_HRxC<I=R_x#HC02RE
CMRCRs0MksRO8_IC;
D
#CRCRs0MksROI_IC;
MH8RVC;
Mo8RCL0_F8FD;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSS8SR_FOEH_OCI0H8EI,R_FOEH_OCI0H8E
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=CRo0F_LF5D8o_C0#CHx50oC_lMk_DOCDI#5HE80,_R8OHEFOIC_HE802C,o0k_MlC_OD5D#80CbE8,R_FOEH_OC80CbE,22
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0oC_x#HCC5o0k_MlC_OD5D#I0H8EI,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,IE_OFCHO_b8C02E2,S
SSSSSSSSSSRRRRH5I8-0E482/_FOEH_OCI0H8E5,RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=o_C0LDFF8C5o0H_#xoC5CM0_kOl_C#DD58IH0RE,8E_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0ERO8_EOFHCC_8b20E2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRRR5b8C04E-2_/8OHEFO8C_CEb0,8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4SOR
F0M#NRM0xFCsR#:R0D8_FOoH_OPC05FsOHEFOIC_HE80*8IH0ME_kOl_C#DD-8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2O;
F0M#NRM0#NsPDD_#PRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#R-48MFI0jFR2=R:RsxCFRR&#H0sM#o.DsP5#80_N20N;F
OMN#0M#0RsDPNR#:R0MsHoE5OFCHO_8IH0IE*HE80_lMk_DOCD8#RF0IMF2R4RR:=#.DP#H0sM#o5sDPN_P#D2-;
-CRLoRHMLODF	NRsllRHblDCCNM00MHFRo#HM#ND
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L.k#RF:RkL0_k_#.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjU,R*8IH0ME_kOl_C#DD+8(RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:URR0Fk_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj4,RnH*I8_0EM_klODCD#6+4RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#nRR:F_k0L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0##2
HNoMDkRF0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05Fs80CbEk_MlC_OD-D#4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNFDRks0_CRo4:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RFOEFR#CLIC0CRCM7RQhNRM8Fbk0kF0RVDRAFRO	)
qv#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C)sRq)77
o#HMRNDI_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoN)DRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7)q7#)
HNoMDqRW7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW7q7)H
#oDMNRh7Q_b0lR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM7CRQ#h
HNoMD RW_b0lR#:R0D8_FOoH;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW- 
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD-#
-CRLoRHM#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCM0_knl_cC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbEc/n;R
RH5VR5b8C0lERFn8Rc>2RR2cURC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mlc_n;k
VMHO0FoMRCD0_CFV0P_Csd8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERFn8Rc
2;CRM8o_C0D0CVFsPC_;d.
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5b8C0;E2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P_Csd8.5CEb02O;
F0M#NRM0M_klODCD_Rd.:MRH0CCos=R:R0oC_lMk_5d.D0CVFsPC_2d.;F
OMN#0MD0RCFV0P_Cs4:nRR0HMCsoCRR:=o_C0D0CVFsPC5VDC0CFPs._d,.Rd2O;
F0M#NRM0M_klODCD_R4n:MRH0CCos=R:R0oC_lMk_54nD0CVFsPC_24n;0

$RbCF_k0L_k#0C$b_#ncRRH#NNss$MR5kOl_C_DDn8cRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bdC_.H#R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_#4nRRH#NNss$MR5kOl_C_DD48nRF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L_k#nRc#:kRF0k_L#$_0bnC_cR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#dR.#:kRF0k_L#$_0bdC_.R#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0L_k#4Rn#:kRF0k_L#$_0b4C_nR#;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRNDI_s0C#M_R#:R0D8_FOoH_OPC05FsM_klODCD_Rnc8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR0Is__CMd:.RR8#0_oDFH
O;#MHoNIDRsC0_Mn_4R#:R0D8_FOoH;H
#oDMNR_HMs_Co#RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soR_#:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C#o_R#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNR8IN_osC_:#RR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFsI_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2-
-R8CMRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDN#
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HMRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRs&RNs8_Cjo52S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRI&RNs8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj"jjRs&RNs8_C4o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRI&RNs8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjj"jjRs&RNs8_C.o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&NRI8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj&"RR8sN_osC58dRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjj"jjRI&RNs8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&s_N8s5CocFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjj&"RR8sN_osC586RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjjRj"&NRI8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj&"RR8sN_osC58nRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjj&"RR8IN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj"jjRs&RNs8_C(o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjjjjjRj"&NRI8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_CUo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj&"RR8IN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_soR5g8MFI0jFR2S;
SIDF_8IN8<sR=jR"j"jjRI&RNs8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co48jRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj&"RR8IN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o54FR8IFM0R;j2
DSSFII_Ns88RR<=""jjRI&RNs8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co48.RF0IMF2Rj;S
SD_FII8N8s=R<R''jRI&RNs8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=NRs8C_sod54RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=NRI8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR7amzRR<=F_k0s5CoI0H8ER-48MFI0jFR2
;
RRRR-Q-RVsR5Ns88_osC2CRso0H#C)sRq)77RHk#MmoRB
piRRRRzs4nRRR:H5VRs8N8sC_soo2RCsMCN
0C-R-RRRRRRsRbF#OC#mR5B,piR7)q7R)2LHCoM-
-RRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CM-R-RRRRRRRRRRRRRRNRs8C_so=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;-
-RRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8sRbF#OC#-;
-MSC8CRoMNCs0zCR4;ns
R--RzRR4R(s:VRHRF5M0NRs8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRs8C_so=R<R7)q7
);S8CMRMoCC0sNC4Rzn
s;
-S-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRmW_B
piRRRRzI4nRRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0CzI4n;R
RR4Rz(:IRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)S;
CRM8oCCMsCN0R(z4I
;
RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
RRzRS4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.j
-S-RRQV58N8s8IH0<ER=cR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.Sz4RR:H5VRNs88I0H8E=R<R24cRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv4Undc7X4RD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5ND[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#"aA7"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*d4nURc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*d4nURc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_ncdUXR47:qR)vnA4__141S4
RRRRRRRRRRRRb0FsRblNRQ57q25jRR=>HsM_C[o52q,R7q7)RR=>D_FII8N8sd54RI8FMR0FjR2,7RQA=">RjR",q)77A>R=RIDF_8sN84s5dFR8IFM0R,j2
SSSSq hRR=>Wh_ ,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R, hR)11A>R=Ra)1, RWA>R=R''j,pRBi=AR>BRmp
i,SRSSR7RRm=qR>bRFCRM,75mAj=2R>kRF0k_L#H45,2[2;R

RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCR
RRzRS.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.Sz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;.6
-S-RRQV58N8s8IH0<ER=dR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRR.SznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.n
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_gU4.7X.RD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5ND.+*[.FR8IFM0R[.*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5UH*42g.R"&RW&"RR0HMCsoC'NHlo[C5*R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42U.4g,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*.;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gU4.7X.R):Rq4vAn._1_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2S,
SRSRRhR q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5R42=F>RkL0_k5#.H*,.[2+4,mR7A25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CRRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSSSSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_cgcnX7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5[c*+8cRF0IMF*Rc[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvcnjgXRc7:NRDLRCDH"#RA"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5Hcnjg2RR&"RW"&MRH0CCosl'HN5oC[2*cR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*gcjn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4c2*2S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSSq7mRR=>FMbC,mR7A25dRR=>F_k0Lck#5RH,c+*[dR2,75mA.=2R>kRF0k_L#Hc5,[c*+,.2RS
SSmS7A254RR=>F_k0Lck#5cH,*4[+27,RmjA52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCR
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
S0SN0LsHkR0CGbO_s#FbRRFVAv)q_c.jU7XURD:RNDLCRRH#"QW)av _m_7 q =)qw7_Qa)1,)R1e_qpAR="&sR#P5NDg+*[gFR8IFM0R[g*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5.H*j2cUR"&RW&"RR0HMCsoC'NHlo[C5*Rg2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42.Ujc,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*g;S
SSoLCHRM
RRRRRRRRRSRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,piRS
SSmS7q>R=RCFbM7,Rm(A52>R=R0Fk_#LkU,5HU+*[(R2,75mAn=2R>kRF0k_L#HU5,[U*+,n2RS
SSmS7A256RR=>F_k0LUk#5UH,*6[+27,RmcA52>R=R0Fk_#LkU,5HU+*[cR2,75mAd=2R>kRF0k_L#HU5,[U*+,d2RS
SSmS7A25.RR=>F_k0LUk#5UH,*.[+27,Rm4A52>R=R0Fk_#LkU,5HU+*[4R2,75mAj=2R>kRF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQu5Rj2=H>RMC_so*5g[2+U,QR7u=AR>jR""R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmRuq=F>Rb,CMRu7mA25jRR=>bHNs0L$_k5#UH2,[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0RC
RSRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM58sN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR") Qa_7vm =_q)7 q_)wQ1Ra,1q)ep=_A"RR&#NsPDU54*4[+UFR8IFM0R*4U[2+4R"&R,)RWQ_a v m7_"A=RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#"aA7"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*.4jc&2RR""WRH&RMo0CCHs'lCNo54[*U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+442*j,.cRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*24U;S
SSoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,piRS
SSmS7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RS
SSmS7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RS
SSmS7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RS
SSmS7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RSSSS75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RS
SSmS7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"Ru7mq>R=RCFbMR,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>NRbs$H0_#Lk4Hn5,[.*+,42Ru7mA25jRR=>bHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_dn1
dnSUzdNRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CSRRRRgzdNRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSzj:NRRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRs_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)v4_6..Xd7RR:DCNLD#RHR)"WQ_a v m7_)q= _q7w1Q)a1,R)peq_"A=R#&RsDPN5*dn[n+dRI8FMR0Fd[n*+R42&,R"RQW)av _m_7 AR="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#AR"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo56H*4R.2&WR""RR&HCM0o'CsHolNC*5[dRn2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*426,4.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*2dn;S
SSoLCHSM
SASS)_qv6X4.dR.7:qR)vnA4_n1d_n1d
RRRRRRRRRRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7q7)RR=>D_FII8N8sR5U8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858URF0IMF2Rj,S
SShS q>R=R W_h1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>hR ,1R1)=AR>1R)aW,R =AR>jR''B,RpRiA=m>RB,pi
SSSSq7mRR=>FMbC,mR7A45d2>R=R0Fk_#LkdH.5,*d.[4+d27,RmdA5j=2R>kRF0k_L#5d.H.,d*d[+j
2,SSSS75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2S,
S7SSm.A5n=2R>kRF0k_L#5d.H.,d*.[+nR2,75mA.R62=F>RkL0_k.#d5dH,.+*[.,62RA7m52.cRR=>F_k0Ldk#.,5Hd[.*+2.c,S
SSmS7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
SSSSA7m52.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7Ag542>R=R0Fk_#LkdH.5,*d.[g+427,Rm4A5U=2R>kRF0k_L#5d.H.,d*4[+U
2,SSSS75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42S,
S7SSm4A5c=2R>kRF0k_L#5d.H.,d*4[+cR2,75mA4Rd2=F>RkL0_k.#d5dH,.+*[4,d2RA7m524.RR=>F_k0Ldk#.,5Hd[.*+24.,S
SSmS7A4542>R=R0Fk_#LkdH.5,*d.[4+427,Rm4A5j=2R>kRF0k_L#5d.H.,d*4[+jR2,75mAg=2R>kRF0k_L#5d.H.,d*g[+2S,
S7SSmUA52>R=R0Fk_#LkdH.5,*d.[2+U,mR7A25(RR=>F_k0Ldk#.,5Hd[.*+,(2RA7m5Rn2=F>RkL0_k.#d5dH,.+*[n
2,SSSS75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2
SSSSA7m5R.2=F>RkL0_k.#d5dH,.+*[.R2,75mA4=2R>kRF0k_L#5d.H.,d*4[+27,RmjA52>R=R0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,QR7u=AR>jR"j"jj,mR7u=qR>bRFC
M,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udA52>R=RsbNH_0$Ldk#.,5Hc+*[dR2,7Amu5R.2=b>RN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Amu5R42=b>RN0sH$k_L#5d.H*,c[2+4,mR7ujA52>R=RsbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
S
SS8CMRMoCC0sNCcRz.
N;SMSC8CRoMNCs0zCRd;gN
MSC8CRoMNCs0zCRd;UN
M
C8sRNO0EHCkO0sMCRFI_s_COEO
	;

-----
-NRp#H0RlCbDl0CMNF0HM#RHRV8CN0kD

--NEsOHO0C0CksRD#CC_O0sRNlF)VRq_vh)R_WHV#
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;F
OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R580CbERR-442/nR2;RRRRRRRRR-RR-RRyF)VRqnv4XR47ODCD#CRMC88C
b0$CkRF0k_L#$_0bHCR#sRNsRN$5lMk_DOCD8#RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LRk#:kRF0k_L#$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05FsM_klODCD#FR8IFM0R;j2RRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;RRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDNRs8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RR-RR-#RkC08RFCRso0H#CWsRq)77
o#HMRNDD_FIs8N8sRR:#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F58dRF0IMF2Rj;RRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHo
;
LHCoMR

R-RR-VRQR8N8s8IH0<ERRNcR#o#HMjR''FR0RkkM#RC8L#H0
RRRRRz4RH:RVNR58I8sHE80R4=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Coj
2;RRRRRRRRD_FII8N8s=R<Rj"jj&"RR8IN_osC5;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=.o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"j"RR&s_N8s5Co4FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"j&"RR8IN_osC584RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co.FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR''RR&I_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR>do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<R8sN_osC58dRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<I=RNs8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRz6RH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR=QR7hR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRCRM8oCCMsCN0R;zn
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzR(R:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRCRM8oCCMsCN0R;zU
R
RR-R-RRQV58sN8ss_CRo2sHCo#s0CR7)q7k)R#oHMRpmBiR
RRgRzRRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBi),Rq)772CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8sRCo<)=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCgRz;R
RR4RzjRR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8sRCo<)=Rq)77;R
RRMRC8CRoMNCs0zCR4
j;RRRRRRRR
RRRRR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoB
piRRRRzR46RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz6R;
RzRR4:nRRRHV50MFR8IN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8IN_osCRR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4n
R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRR4z4RV:RFHsRRRHMM_klODCD#FR8IFM0RojRCsMCN
0CRRRRRRRR-Q-RVNR58I8sHE80Rc>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z4RH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
.;RRRRRRRR-Q-RVNR58I8sHE80RR<=cM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4d:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR4
d;RRRR-t-RMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4c:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qRD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*24nR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55+*424Rn,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqRv:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDIN_I858sjR2,q=4R>FRDIN_I858s4R2,q=.R>FRDIN_I858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s25d,uR7)Rqj=D>RFsI_Ns885,j2R)7uq=4R>FRDIN_s858s4R2,
RRRRRRRRRRRRRRRRRRRRRRRR7RRu.)qRR=>D_FIs8N8s25.,uR7)Rqd=D>RFsI_Ns885,d2RRW =I>RsC0_M25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRpWBi>R=RiBp,uR7m>R=R0Fk_#Lk5[H,2
2;RRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0Rcz4;R
RRRRRRMRC8CRoMNCs0zCR4
4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0s#CRCODC0N_sl
;

