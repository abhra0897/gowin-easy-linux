--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lbj6j#/L0lbNbC/s#GHHDMDG/HoL/CPM_HCs0Gl/#k3D0PyE84
Rf-
-
---
-HR1o8MCRDvk0DHbHRCsIEH0RbbHCVLk#HR5MNRO#FCRVHRbbHCDMoHM2-
-RsaNoRC0:HRXDGHM

--
LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
H
DLssN$$R#MHbDV
$;kR#C#b$MD$HV30N0skHL03C#N;DD
M
C0$H0RswH#s0uFO8k0H#R#o
SCsMCH
O5SHSI8q0ERH:RMo0CC
s;SHSI8A0ERH:RMo0CCSs
2S;
b0FsRS5
SRqR:MRHR0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2S;
SRAR:MRHR0R#8F_Do_HOP0COFIs5HE80AR-48MFI0jFR2S;
SRqA:kRF00R#8F_Do_HOP0COFIs5HE80AH*I8q0E-84RF0IMF2Rj
-SS-RRA*
RqS
2;CRM8w#Hs0Fus80kO#
;
NEsOHO0C0CksRONsEF4RVHRwsu#0skF8OR0#H
#
R#RRHNoMD_RNNRkG:0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2R;
RHR#oDMNRNL_k:GRR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;C
Lo
HMSsVFNqM8:FRVsNRHRRHMjFR0R8IH0-Eq.CRoMNCs0SC
SsVFNAM8:FRVsLRHRRHMjFR0R8IH0-EA.CRoMNCs0SC
SASq58IH0*EAH+NRR2HLRR<=NN5H2MRN85RLH;L2
CSSMo8RCsMCNR0CVNFsM;8A
HSSVJ_C:VRHRN5HRj=R2CRoMNCs0SC
SASq58IH0-EA4<2R=5RNjN2RML8R58IH0-EA4
2;SMSC8CRoMNCs0HCRVJ_C;S
SHMV_CRJ:H5VRH/NR=2RjRMoCC0sNCS
SS5qAI0H8EHA*NH+I8A0E-R42<5=RMRF0NN5H2N2RML8R58IH0-EA4
2;SMSC8CRoMNCs0HCRVC_MJS;
CRM8oCCMsCN0RsVFNqM8;V
SFMsN8RA:VRFsHHLRMRRj0IFRHE80AR-.oCCMsCN0
qSSAH5I8A0E*H5I8q0E-R42+LRH2=R<RIN5HE80q2-4R8NMRF5M05RLH2L2;C
SMo8RCsMCNR0CVNFsM;8A
qSSAH5I8A0E*H5I8q0E-R42+HRI8A0E-R42<N=R58IH0-Eq4N2RML8R58IH0-EA4
2;CRM8NEsO4
;

LDHs$NsR Q  D;
HNLss#$R$DMbH;V$
Ck#RM#$bVDH$03N0LsHk#0C3DND;#
kC RQ 1 3ap7_mBtQ_n44cD3NDb;
NNO	oeCRBumvmhh aH1R#F
OlMbFCRM0u QuA
zwSsbF0
R5SRSm:kRF00R#8F_Do;HO
QSSRH:RM0R#8F_Do
HOS
2;CRM8ObFlFMMC0
;
Ns00H0LkC$R#MD_LN_O	LRFGFuVRQAu z:wRRlOFbCFMMH0R#sR0k
C;-C-RMF8RVHRbbkCLV-

-MR 8NRLON	IsO8RFNlb0HHLD$H0RlOFbCFMM
0#CRM8evBmu mhh;a1
D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
Ck#RFPOlMbFC#M03DND;C

M00H$8RN8osCR
H#SMoCCOsH5S
SI0H8E:RRR0HMCsoC;S
SI0H8E:qRR0HMCsoC;S
SHCM8G:RRR0HMCsoC;S
SMLklC:sRR0HMCsoC;S
SsRCoR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPD2
S;b
SFRs05S
SBRHM:MRHR8#0_oDFH
O;SRSqRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
SRARRH:RM0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SsRC#:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj
;S2
0SN0LsHkR0C\N3sMR	\:MRH0CCosR;
RNRR0H0sLCk0Rs\3CPlFCF_M_sINM:\RR0HMCsoC;M
C88RN8osC;N

sHOE00COkRsCNEsO4VRFR8N8sRCoHR#
RHR#oDMNR#sCkRD0:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;C
Lo
HMS#sCkRD0<q=RRA+RRO+RH
M;S_HVjH:RVHR5MG8CR4>R2CRoMNCs0
CRSFSVsFDFbRj:VRFsHMRHR0jRFHRI8q0E-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#s;Co
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCRo#:NRDLRCDH4#R;S
SLHCoMS
SSosC#b:RHLbCkSV
SbSSFRs0l5Nb
SSSSQSSRR=>skC#DH052S,
SSSSS=mR>CRs#25H
SSSS
2;SMSC8CRoMNCs0VCRFFsDF;bj
MSC8CRoMNCs0RCRHjV_;S

H4V_:VRHRM5H8RCG=2R4RMoCC0sNCSR
SsVFDbFF.V:RFHsRRRHMjFR0R8IH0-Eq4CRoMNCs0SC
S0SN0LsHkR0C\N3sMR	\FsVRCqo#RD:RNDLCRRH#s;Co
SSSNs00H0LkC3R\sFClPMC_FN_IsRM\FsVRCqo#RD:RNDLCRRH#4S;
SoLCHSM
SCSso:#qRbbHCVLk
SSSSsbF0NRlbS5
SSSSS=QR>CRs#0kD5,H2
SSSSmSSRR=>s5C#HS2
S2SS;S
SCRM8oCCMsCN0RsVFDbFF.S;
CRM8oCCMsCN0RVRH_
4;
VSH_R.:H5VR.M*H8RCG=kRMlsLC2CRoMNCs0
CRSFSVsFDFbRd:VRFsHMRHR8IH0REq0IFRHE80-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHRosC;S
SS0N0skHL0\CR3lsCF_PCMIF_N\sMRRFVs#CoARR:DCNLD#RHR
4;SCSLo
HMSsSSCAo#:HRbbkCLVS
SSFSbsl0RN
b5SSSSSRSQ=s>RCD#k025H,S
SSSSSm>R=R#sC5
H2SSSS2S;
S8CMRMoCC0sNCFRVsFDFb
d;S8CMRMoCC0sNCHRRV;_.
H
SV:_dRRHV5H.*MG8CRM<RkClLso2RCsMCNR0C
VSSFFsDF:bcRsVFRHHRMHRI8q0ERR0FI0H8ER-4oCCMsCN0
SSSNs00H0LkC3R\s	NM\VRFRosC#:BRRLDNCHDR#CRsoS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:BRRLDNCHDR#;R4
LSSCMoH
SSSs#CoBb:RHLbCkSV
SbSSFRs0l5Nb
SSSSQSSRR=>skC#DH052S,
SSSSS=mR>CRs#25H
SSSS
2;SMSC8CRoMNCs0VCRFFsDF;bc
MSC8CRoMNCs0RCRHdV_;M
C8sRNO;E4
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
#
kCORPFFlbM0CM#D3ND
;
CHM00V$RDsFFR
H#SCSoMHCsO
R5SSSSI0H8ERQhRH:RMo0CC:sR=jRg;S
SSHSI8m0Ez:aRR0HMCsoCRR:=6
c;SSSSMLklCRsRRH:RMo0CC:sR=;R6
SSSS8IH0REqRRR:HCM0oRCs:6=R;S
SSMSH8RCGRRRR:MRH0CCos=R:4S
S2S;
SsbF0
R5SSSSQkMb0:RRRMRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2S;
SmSSkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2S
S2S;
S0N0skHL0\CR3MsN	:\RR0HMCsoC;S
SNs00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
MV8RDsFF;N

sHOE00COkRsCNEsO4VRFRFVDFHsR#RR
RORRFFlbM0CMR8N8s
CoSoRRCsMCH5OR
RSRSHSI8R0ERH:RMo0CC
s;SSRRS8IH0REq:MRH0CCosS;
RSRSHCM8G:RRR0HMCsoC;R
SRMSSkClLsRR:HCM0o;Cs
SSSsRCoR:RRR0HMCsoCRR--hCNlRRFV0RECDCCPDR
SR
2;SbRRFRs05S
SBRHM:MRHR8#0_oDFH
O;SRSqRRR:H#MR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;SRSARRR:H#MR0D8_FOoH_OPC05FsR8IH04E-RI8FMR0Fj
2;SCSs#RR:FRk0#_08DHFoOC_POs0F58IH04E-RI8FMR0FjS2
R;R2
RRRCRM8ObFlFMMC0
;
Sb0$CER#H_V00DNLC#RHRsNsN5$RMLklC.s/RI8FMR0FjF2RVMRH0CCos
;
SMVkOF0HMER#HxV0C5sFHCM8GRR:HCM0o2CsR0sCkRsM#VEH0N_0LRDCHS#
SsPNHDNLC0R#C:bRR0HMCsoC;S
SPHNsNCLDRL0NDPC_NRsR:ER#H_V00DNLCS;
LHCoMS
S#b0CRR:=4S;
SsVFRHHRMRR40HFRMG8C-D4RF
FbS#SS0RCb:#=R0RCb*;R.
CSSMD8RF;Fb
VSSFHsRRRHMjFR0RlMkL/Cs.FRDFSb
SNS0L_DCP5NsH:2R=0R#C*bRR*5.H2+4;S
SCRM8DbFF;S
SskC0s0MRNCLD_sPN;C
SM#8RE0HVxFCs;S

O#FM00NMRMDCoRE0:MRH0CCos=R:R8IH0MEQ/lMkL;Cs
FSOMN#0MI0RHE80ARR:HCM0oRCs:D=RCEMo0RR-I0H8E
q;
FSOMN#0M#0RE0HVNC88sRR:#VEH0N_0LRDC:#=RE0HVxFCs58HMC;G2
C
Lo
HMSsVFDbFF_R4:VRFs[MRHR04RFkRMlsLC/o.RCsMCN
0CSoLCHSM
RsRRCqo#:8RN8osC
RSRRMoCCOsHRblNRS5
S8IH0=ER>CRDM0oE-H#EV80N85Cs[2-4-
4,SHSI8q0ERR=>I0H8E
q,SMSH8RCG=[>R,S
SMLklC=sR>kRMlsLC,S
SsRCoR>R=R8HMCSG
R2RR
RSRRsbF0NRlbS5
RSRRRHRBM>R=RbQMkD05CEMo0.*5*4[-2R2,
RSRRRRRq>R=RbQMkD05CEMo0.*5*4[-2R-48MFI0DFRCEMo0**.54[-2E+#HNV08s8C54[-22+4,R
SRRRRR=AR>MRQb5k0DoCME.0**4[-RI8FMR0FDoCME50*.-*[4#2+E0HVNC88s-5[442+2S,
RRRRRCRs#>R=R0mkb5k0DoCME[0*-84RF0IMFCRDM0oE*-5[4#2+E0HVNC88s-5[442+2R
SR;R2
RSRRR--OsNs$FRVsER0CCRMGV0RDsFF
VSSFFsDFjb_:FRVsRRHHjMRRR0F#VEH08N8C[s5--42#VEH08N8Cjs52CRoMNCs0RC
RRRSRSRSmbk0kD05CEMo0[*5-+42RRH2<'=Rj
';SMSC8CRoMNCs0VCRFFsDFjb_;S

R-RR-DRNs8CN$CRoMNCs0
C8SFSVsFDFb:_NRsVFRHHRMRRj0#FRE0HVNC88s25j-o4RCsMCN
0CSNSS0H0sLCk0Rs\3N\M	RRFVs#CoRD:RNDLCRRH#HCM8GS;
S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#RR:DCNLD#RHR
4;SCSLo
HMSsSSC:o#RbbHCVLk
SSSSFSbsl0RN
b5SSSSSQSSRR=>QkMb0C5DM0oE*5.*[2-4+H#EV80N85Cs[2-4-H#EV80N85Csj42++,H2
SSSSSSSm>R=R0mkb5k0DoCME50*[2-4+#H+E0HVNC88s-5[4#2-E0HVNC88s25j+
42SSSSS2SS;S
SCRM8oCCMsCN0RsVFDbFF_
N;
MSC8CRoMNCs0VCRFFsDF4b_;S

H#V_FNk#:VRHRk5MlsLCR8lFR=.RRR42oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVsOCoN$ss#RR:DCNLD#RHR8HMC
G;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosCOsNs$:#RRLDNCHDR#;R4
CSLo
HMSRRRVDFsF_FbdV:RFHsRRRHM4FR0RCRDM0oE-H#EV80N85CsMLklC.s/2+-4#VEH08N8Cjs52CRoMNCs0SC
S0N0skHL0\CR3MsN	F\RVCRso:#RRLDNCHDR#MRH8;CG
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRso:#RRLDNCHDR#;R4
RSRRoLCHSM
RRRRRCRsoR#:bCHbL
kVSRRRRbRRFRs0l5Nb
RSRRRRRRQRRRR=>QkMb0H5I8Q0Eh2-H,R
SRRRRRRRRm>R=R0mkb5k0I0H8Eamz-
H2SRRRR2RR;R
SRMRC8CRoMNCs0VCRFFsDFdb_;R
SRCRsosONs:$#RbbHCVLk
RSRRRRRb0FsRblN5R
SRRRRRRRRQ>R=RbQMkI05HE80QDh-CEMo0
2,SRRRRRRRRRRm=m>Rkk0b0H5I8m0EzDa-CEMo0S2
RRRRR;R2
RSRR0mkb5k0I0H8Eamz-MDCo+E0#VEH08N8CMs5kClLs2/.-H#EV80N85Csj82RF0IMFHRI8m0EzDa-CEMo02+4RR<=
SSSSMSQb5k0I0H8E-QhDoCME#0+E0HVNC88sk5MlsLC/-.2#VEH08N8Cjs52FR8IFM0R8IH0hEQ-MDCo+E04R2;
MSC8CRoMNCs0HCRVF_#k;#N
8CMRONsE
4;



DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00V$RDsFF_8N8CHsR#S
SoCCMsRHO5S
SSHSI8Q0Eh:RRR0HMCsoCRR:=g
j;SSSSI0H8EamzRH:RMo0CC:sR=cR6;S
SSkSMlsLCR:RRR0HMCsoCRR:=6S
S2S;
SsbF0
R5SSSSQkMb0:RRRMRHR8#0_oDFHPO_CFO0sH5I8Q0EhR-48MFI0jFR2S;
SmSSkk0b0RR:FRk0#_08DHFoOC_POs0F58IH0zEmaR-48MFI0jFR2S
S2C;
MV8RDsFF_8N8C
s;
ONsECH0Os0kCsRNORE4FVVRDsFF_8N8CHsR#SR
O#FM00NMRMDCoRE0:MRH0CCos=R:R8IH0MEQ/lMkL;Cs
oLCHSM
VDFsF_Fb4V:RF[sRRRHM4FR0RlMkL/Cs.CRoMNCs0SC
S0mkb5k0DoCME[0*-84RF0IMFCRDM0oE*-5[442+2=R<RMRQb5k0DoCME50*.-*[442-RI8FMR0FDoCME.0**-5[442+2S
SSSSSSSSSSRSRRQ+RM0bk5MDCo*E0.-*[4FR8IFM0RMDCo*E05[.*-+424S2
SSSSSSSSSRSSRRR+QkMb0C5DM0oE**5.[2-42
;
SkSm00bk5MDCo*E054[-2<2R=jR''S;
CRM8oCCMsCN0RsVFDbFF_
4;
VSH_k#F#RN:H5VRMLklClsRF.8RR4=R2CRoMNCs0SC
S0mkb5k0I0H8Eamz-84RF0IMFHRI8m0EzDa-CEMo0<2R=MRQb5k0I0H8E-Qh4FR8IFM0R8IH0hEQ-MDCo2E0;SR
CRM8oCCMsCN0R_HV##FkN
;
CRM8NEsO4
;
DsHLNRs$HCCC;kR
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3ND
;
CHM00N$R8s8CaCsC.#RH
CSoMHCsOS5
S8IH0REq:MRH0CCosS;
S8IH0REA:MRH0CCosS;
SC0sCRRR:MRH0CCos2
S;b
SFRs05S
Sqq,RlA,RRH:RM0R#8F_Do;HO
qSSA:RRRRHM#_08DHFoOC_POs0F58IH0*EAI0H8E4q-RI8FMR0Fj
2;SsSbFO8k0RR:FRk0#_08DHFoOC_POs0F58IH0+EAI0H8E4q-RI8FMR0FjS2
SR--ARR*q2
S;M
C88RN8aCss.CC;

RNEsOHO0C0CksRONsEF4RV8RN8aCss.CCR
H#RORRF0M#NRM00EECHRoE:0R#8F_Do_HOP0COF4s56FR8IFM0RRj2:B=Rm_he1_a7pQmtB _eB)am58IH0-Eq44,Rn
2;RORRFFlbM0CMRFVDFRs
RRRRRMoCCOsHRS5
SHSI8Q0Eh:RRR0HMCsoCRS;
SHSI8m0Ez:aRR0HMCsoCRS;
SkSMlsLCR:RRR0HMCsoCRS;
SHSI8q0ER:RRR0HMCsoCRS;
SMSH8RCGR:RRR0HMCsoC
RRRR2RR;R
RRRRRRsbF0
R5RRRRRRRRRRRRRMRQbRk0RH:RM0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;RRRRRRRRRRRRRkRm00bkRF:Rk#0R0D8_FOoH_OPC05FsI0H8Eamz-84RF0IMF2Rj
RRRRRRR2R;
RMRC8FROlMbFC;M0
R
RRlOFbCFMMV0RDsFF_8N8CRs
RRRRRMoCCOsHRS5
SHSI8Q0Eh:RRR0HMCsoCRS;
SHSI8m0Ez:aRR0HMCsoCRS;
SkSMlsLCR:RRR0HMCsoC
RRRR2RR;R
RRRRRRsbF0
R5RRRRRRRRRRRRRMRQbRk0RH:RM0R#8F_Do_HOP0COFIs5HE80Q4h-RI8FMR0Fj
2;RRRRRRRRRRRRRkRm00bkRF:Rk#0R0D8_FOoH_OPC05FsI0H8Eamz-84RF0IMF2Rj
RRRRRRR2R;
RMRC8FROlMbFC;M0
R
RRMVkOF0HMCR8bW0EHE80R0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRsVFRHHRM6R4RI8FMR0FjFRDFSb
H5VR0EECH5oEH=2RR''42ER0CSM
RsRRCs0kM+RH4S;
CRM8H
V;RRRRR8CMRFDFbR;
RRRRskC0sjMR;R
RR8CMRb8C0HEW8;0E
R
RRMOF#M0N0CR8bR0E:MRH0CCos=R:Rb8C0HEW8;0E
RRRO#FM00NMR8IH0RE0:MRH0CCos=R:R8IH0+EAI0H8E.q+;R
RRb0$CHRDlH#R#sRNsRN$5b8C04E+RI8FMR0FjF2RVMRH0CCosR;

RRRVOkM0MHFRDONOlhkL#CsR0sCkRsMD#HlR
H#RRRRRNRPsLHND0CREMC_kClLs:#RRlDH#R;
RCRLo
HMRRRRRER0Ck_MlsLC#25jRR:=I0H8E
q;RRRRRFRVsRRHH4MRRR0F80CbER+4DbFF
RRRRRRRRER0Ck_MlsLC#25HRR:=0_ECMLklC5s#H2-4/+.RRE50Ck_MlsLC#-5H4l2RF.8R2R;
RRRRR8CMRFDFbR;
RRRRR0sCkRsM0_ECMLklC;s#
RRRR8CMRDONOlhkL#Cs;

RRORRF0M#NRM0MLklCRs#:HRDl:#R=NRODkOhlsLC#R;

RRRVOkM0MHFRDONOlpHR0sCkRsMD#HlR
H#RRRRRNRPsLHND0CREDC_HRl#:HRDl
#;RRRRRNRPsLHNDMCRkRlL:MRH0CCosR;
RCRLo
HMRRRRRER0CH_Dlj#52=R:R
j;RRRRRkRMl:LR=HRI8q0E;R
RRRRRVRFsHMRHR04RFCR8b+0E4FRDFRb
SC0E_lDH#25HRR:=0_ECD#Hl54H-2RR+MLkl*8IH0;E0
MRSkRlL:M=Rk/lL.RR+5lMkLFRl82R.;R
RRRRRCRM8DbFF;R
RRRRRskC0s0MREDC_H;l#
RRRR8CMRDONOlpH;

RRORRF0M#NRM0PDCOH:lRRlDH#=R:RDONOlpH;R
RRo#HMRNDL0HosRCC:0R#8F_Do_HOP0COFPs5CHODlC58b+0E442-RI8FMR0Fj
2;R#RRHNoMDNROs,s$Ro#HM#,RH4oMR#:R0D8_FOoH;L

CMoHRH
SVC_	CNb_8s8CaCsC:VRHRs50C=CRRRj2oCCMsCN0RR--kR#CVRFsbCHbDHHMMNoRMD8RFOIRF
#0
#SSHRoM<q=RRsGFR
A;SHS#oRM4<q=RRRFsAS;
SsONs<$R=MR5Fq0RlN2RMA8R;S
SL0Hos5CCI0H8E40-RI8FMR0Fj<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E
q2SSSSSSSSSRS&OsNs$S
SSSSSSSSS&ARq58IH0-EA4FR8IFM0R
j2SSSSSSSSSRS&Bemh_71a_tpmQeB_ mBa),5jR;42
S
SVNFsM:8qRsVFRRHNH4MRRR0FI0H8Edq-RMoCC0sNCS
SSoLH0CsC5N5H+*42I0H8E40-RI8FMR0FHIN*HE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,I0H8E4q+-2HN
SSSSSSSSSSSS&SSR5qAI0H8E5A*H4N+2R-48MFI0IFRHE80AN*H2S
SSSSSSSSSSSSS&mRBh1e_ap7_mBtQ_Be a5m)jH,RN2+4;S
SCRM8oCCMsCN0RsVFNqM8;S
S-F-RMLCRCsVFCER0CNRD#P0RCFO0sS
SL0Hos5CC58IH0-Eq4I2*HE800R-48MFI05FRI0H8E.q-2H*I800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)j.,R2S
SSSSSSSSSSSSSSRS&#MHo
SSSSSSSSSSSSSSSSq&RAH5I8A0E*H5I8q0E--424FR8IFM0R8IH0*EA58IH0-Eq.
22SSSSSSSSSSSSSSSS&mRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q2-4;S
S-D-RNR#0P0COFSs
SoLH0CsC58IH0*EqI0H8E40-RI8FMR0F58IH0-Eq4I2*HE800<2R=SR
SSSSSSSSSSSSSBSSm_he1_a7pQmtB _eB)am5Rj,4S2
SSSSSSSSSSSSSRS&#MHo4S
SSSSSSSSSSSSSSq&RAH5I8A0E*8IH0-Eq4FR8IFM0R8IH0*EA58IH0-Eq4
22SSSSSSSSSSSSS&SSRhBmea_17m_pt_QBea Bmj)5,HRI8q0E-
42SSSSSSSSSSSSS&SSR
q;
VSSFFsDF:b.VRFs[MRHR04RFCR8bR0EoCCMsCN0
SSSlR4:RFVDFSs
SoSSCsMCHlORN5bR
SSSSSSSI0H8ERQhRR=>PDCOH[l52RR-PDCOH[l5-,42
SSSSSSSI0H8EamzRR=>PDCOH[l5+R42-CRPOlDH5,[2
SSSSSSSMLklCRsRRR=>MLklC5s#[2-4,S
SSSSSS8IH0REqR>R=R8IH0,Eq
SSSSSSSHCM8GRRRRR=>[S
SS
S2SSSSb0FsRblNRS5
SSSSSMSQbRk0R=RR>HRLoC0sCC5POlDH5-[24FR8IFM0ROPCD5Hl[2-42S,
SSSSSkSm00bkR=RR>HRLoC0sCC5POlDH54[+2R-48MFI0PFRCHODl25[2S
SS;S2
CSSMR8RoCCMsCN0RsVFDbFF.S;
CRM8oCCMsCN0R_HV	bCC_8N8CssaC
C;
VSH_0MF	bCC_8N8CssaCRC:H5VR0CsCR4=R2CRoMNCs0-CR-#RkCVRHR8N8CNsRVs0CRC0ERDlk0DHbH
CsS-S-R8IH0REq>c=R
#SSHRoMRR<=qFRGs;RA
#SSH4oMRR<=qsRFR
A;SNSOsRs$<5=RMRF0qRl2NRM8AS;
SoLH0CsC58IH0-E04FR8IFM0RRj2<R=RBemh_71a_tpmQeB_ mBa),5jR8IH02Eq
SSSSSSSS&SSRsONsS$
SSSSSSSSSq&RAH5I8A0E-84RF0IMF2Rj
SSSSSSSS&SSRhBmea_17m_pt_QBea Bmj)5,2R4;S

S_HVI0H8ERq:H5VRI0H8E>qRRRd2oCCMsCN0
SSSL0Hos5CC.H*I800E-84RF0IMFHRI800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)jI,RHE80qS2
SSSSSSSSSSSS&ARq5I.*HE80AR-48MFI0IFRHE80AS2
SSSSSSSSSSSS&
RqSSSSSSSSSSSSSq&R;S

SFSVs8NMqV:RFHsRNMRHR0.RFHRI8q0E-odRCsMCN
0CSSSSL0Hos5CC5+HN4I2*HE800R-48MFI0HFRNH*I800E2=R<RmRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q-+4H
N2SSSSSSSSSSSSS&SSR5qAI0H8E5A*H4N+2R-48MFI0IFRHE80AN*H2S
SSSSSSSSSSSSSSq&R
SSSSSSSSSSSSSSS&mRBh1e_ap7_mBtQ_Be a5m)jH,RN
2;SCSSMo8RCsMCNR0CVNFsM;8q
SSS-F-RMLCRCsVFCER0CNRD#P0RCFO0sS
SSoLH0CsC5H5I8q0E-*42I0H8E40-RI8FMR0F58IH0-Eq.I2*HE800<2R=BRRm_he1_a7pQmtB _eB)am5Rj,.S2
SSSSSSSSSSSSSSSS&HR#oSM
SSSSSSSSSSSSSSSS&ARq58IH0*EA58IH0-Eq442-RI8FMR0FI0H8E5A*I0H8E.q-2S2
SSSSSSSSSSSSSSSS&
RqSSSSSSSSSSSSSSSSSB&Rm_he1_a7pQmtB _eB)am5Rj,I0H8E.q-2S;
S8CMRMoCC0sNCVRH_8IH0;Eq
S
SHIV_HE80q:_jRRHV58IH0REq=2RdRMoCC0sNCS
SSR--FRMCLFCVs0CREDCRNR#0P0COFSs
SHSLoC0sC*5.I0H8E40-RI8FMR0FI0H8ER02<R=RBemh_71a_tpmQeB_ mBa),5jR
.2SSSSSSSSSSSSS#&RH
oMSSSSSSSSSSSSSq&RA*5.I0H8E4A-RI8FMR0FI0H8E
A2SSSSSSSSSSSSSq&R
SSSSSSSSSSSSRS&q
;
SMSC8CRoMNCs0HCRVH_I8q0E_
j;S-S-R#DN0CRPOs0F
LSSHso0CIC5HE80qH*I800E-84RF0IMFIR5HE80q2-4*8IH02E0RR<=RhBmea_17m_pt_QBea Bmj)5,2R4
SSSSSSSSSSSSSSS&HR#o
M4SSSSSSSSSSSSS&SSR5qAI0H8EIA*HE80qR-48MFI0IFRHE80AI*5HE80q2-42S
SSSSSSSSSSSSSSq&R
SSSSSSSSSSSSSSS&mRBh1e_ap7_mBtQ_Be a5m)jI,RHE80q2-4;S

SsVFDbFFdF:VsRR[H4MRRR0F80CbECRoMNCs0SC
S4Sl:VRRDsFF_8N8CSs
SoSSCsMCHlORN5bR
SSSSSSSI0H8ERQhRR=>PDCOH[l52RR-PDCOH[l5-,42
SSSSSSSI0H8EamzRR=>PDCOH[l5+R42-CRPOlDH5,[2
SSSSSSSMLklCRsRRR=>MLklC5s#[2-4
SSSSS2
SbSSFRs0lRNb5S
SSSSSSbQMkR0RR>R=RoLH0CsC5OPCD5Hl[42-RI8FMR0FPDCOH[l5-242,S
SSSSSS0mkbRk0R>R=RoLH0CsC5OPCD5Hl[2+4-84RF0IMFCRPOlDH52[2
SSSS
2;SMSC8oRRCsMCNR0CVDFsFdFb;C
SMo8RCsMCNR0CHMV_FC0	CNb_8s8CaCsC;S

b8sFkRO0<L=RHso0CPC5CHODlC58b+0E4.2-RI8FMR0FPDCOH8l5CEb022+4;
R
CRM8NEsO4
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;
LDHs$NsRM#$bVDH$k;
##CR$DMbH3V$Ns00H0LkCN#3D
D;
Ck#RFPOlMbFC#M03DND;R
RRRRR
0CMHR0$#DlNDDvk0#RH
CSoMHCsOS5
SHNI8R0E:MRH0CCos=R:R
g;SISLHE80RH:RMo0CC:sR=;Rg
ISSHE80RRR:HCM0oRCs:4=RU2
S;b
SFRs05S
SqRRRRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;SRSAR:RRRRHMR8#0_oDFHPO_CFO0sI5LHE80-84RF0IMF2Rj;S
Su7)mRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S
S-A-RRq*R
;S2
0SN0LsHkR0C\N3sMR	\:MRH0CCosS;
Ns00H0LkC3R\sFClPMC_FN_IsRM\:MRH0CCosC;
M#8RlDNDv0kD;N

sHOE00COkRsCNEsO4VRFRN#lDkDvDH0R#R

RkRVMHO0F#MRkIb5HE80NI,RHE80LRR:HCM0o2CsR0sCkRsMHCM0oRCsHR#
RCRLo
HMRRRRRVRHRH5I8N0ERI>RHE80L02RE
CMSCRs0MksR8IH0;EN
RRRRCRRD
#CRsSRCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRM#8Rk
b;
RRRVOkM0MHFRVHM58IH0,ENR8IH0REL:MRH0CCoss2RCs0kMMRH0CCos#RH
RRRLHCoMR
RRRRRH5VRI0H8E<NRR8IH02ELRC0EMR
SskC0sIMRHE80NR;
RRRRR#CDCs
SCs0kMHRI8L0E;R
RRRRRCRM8H
V;RCRRMH8RM
V;
RRRO#FM00NMR8IH0REq:MRH0CCos=R:RVHM5HNI8,0ERHLI820E;R
RRMOF#M0N0HRI8A0ERH:RMo0CC:sR=kR#bI5NHE80,IRLHE802
;
RORRFFlbM0CMRswH#s0uFO8k0S#
oCCMs5HO
ISSHE80qRR:HCM0o;Cs
ISSHE80ARR:HCM0o
CsS
2;SsbF0
R5SRSqRH:RM#RR0D8_FOoH_OPC05FsN8IH04E-RI8FMR0Fj
2;SRSARH:RM#RR0D8_FOoH_OPC05FsL8IH04E-RI8FMR0Fj
2;SASqRF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2S
S-A-RRq*R
;S2
RRRCRM8ObFlFMMC0
;
RORRFFlbM0CMR8N8CssaC
C.SMoCCOsH5S
SI0H8E:qRR0HMCsoC;S
SI0H8E:ARR0HMCsoC;S
S0CsCR:RRR0HMCsoC
;S2
FSbs50R
qSS,lRq,RRA:MRHR8#0_oDFH
O;SASqRRR:H#MR0D8_FOoH_OPC05FsL8IH0NE*I0H8ER-48MFI0jFR2S;
SFbs80kORF:Rk#0R0D8_FOoH_OPC05FsL8IH0NE+I0H8ER-48MFI0jFR2S
S-A-RRq*R
;S2
RRRCRM8ObFlFMMC0
;
R#RRHNoMD_RNNRkG:0R#8F_Do_HOP0COFIs5HE80qR-48MFI0jFR2R;
RHR#oDMNRNL_k:GRR8#0_oDFHPO_CFO0sH5I8A0E-84RF0IMF2Rj;R
RRo#HMRNDNRLRRRR:#_08DHFoOC_POs0F5HNI8*0EL8IH04E-RI8FMR0Fj
2;R#RRHNoMDCRs#0kD:0R#8F_Do_HOP0COFNs5I0H8EI+LHE80-84RF0IMF2Rj;C
LoRHM
RRR-1-RIRNbqMRN8RRAHMVRC#OC#$Ns
RRRHDVqNCsosRA:H5VRN8IH0>ERRHLI820ERMoCC0sNCR
RRRRRVDFsF.Fb:FRVsRRHHjMRRR0FL8IH04E-RMoCC0sNCS
SNs00H0LkC3R\s	NM\VRFRosC#:qRRLDNCHDR#;Rj
NSS0H0sLCk0Rs\3CPlFCF_M_sINMF\RVCRsoR#q:NRDLRCDH4#R;R
RRNSS0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RSRRosC#Rq:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RAH
2,SRRRRmRRRR=>Nk_NG25H
RSRR
2;SRRRs#CoAb:RHLbCkSV
RbRRFRs0l5Nb
RSRRRRRQ>R=RHq52S,
RRRRRRRm=L>R_GNk5
H2SRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
.;RRRRRFRVsFDFbR4:VRFsHMRHRHLI8R0E0NFRI0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#CoARR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:ARRLDNCHDR#;R4
RRRRLRRCMoH
RSRRosC#RA:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RqH
2,SRRRRmRRRR=>Lk_NG25H
RSRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;b4
RRRCRM8oCCMsCN0RqHVDoNsC;sA
R
RRqHV#DlNDACs:VRHRI5NHE80RR<=L8IH0RE2oCCMsCN0
RRRRVRRFFsDF:bNRsVFRHHRMRRj0NFRI0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#CoBRR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:BRRLDNCHDR#;R4
NSS0H0sLCk0Rs\3N\M	RRFVs#Co1RR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:1RRLDNCHDR#;R4
RRRRLRRCMoH
RSRRosC#RB:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RqH
2,SRRRRmRRRR=>Nk_NG25H
RSRR
2;SRRRs#Co1b:RHLbCkSV
RbRRFRs0l5Nb
RSRRRRRQ>R=RHA52S,
RRRRRRRm=L>R_GNk5
H2SRRR2R;
RRRRR8CMRMoCC0sNCFRVsFDFb
N;RRRRRFRVsFDFbRL:VRFsHMRHRHNI8R0E0LFRI0H8ER-4oCCMsCN0
NSS0H0sLCk0Rs\3N\M	RRFVs#Co7RR:DCNLD#RHR
j;S0SN0LsHkR0C\C3slCFP__MFIMNs\VRFRosC#:7RRLDNCHDR#;R4
RRRRLRRCMoH
RSRRosC#R7:bCHbL
kVSRRRb0FsRblN5R
SRRRRR=QR>5RAH
2,SRRRRmRRRR=>Lk_NG25H
RSRR
2;RRRRRMRC8CRoMNCs0VCRFFsDF;bL
RRRCRM8oCCMsCN0RqHV#DlNDACs;R

RHRws1#00:CbRswH#s0uFO8k0S#
oCCMsRHOlRNb5S
SI0H8E=qR>HRI8q0E,S
SI0H8E=AR>HRI8A0E

S2SsbF0NRlb
R5SRSq=N>R_GNk,S
SA>R=RNL_k
G,SASqRR=>NSL
2
;
RqRR8s8CaCsC.:HRR8N8CssaC
C.SMoCCOsHRblNRS5
S8IH0REq=I>RHE80qS,
S8IH0REA=I>RHE80AS,
SC0sCRRR=j>RS-SS-RR4HNVR8s8CR0NVC0sRElCRkHD0bCDHsj,RR#CDC2
S
FSbsl0RN5bR
qSSl>R=RNN_kjG52S,
SRqR=N>R_GNk58IH0-Eq4
2,SRSARR=>Lk_NGH5I8A0E-,42
qSSA>R=R,NL
bSSskF8O=0R>CRs#0kD
;S2
H
SVF_I:VRHRH5I8R0E<I=RHE80qRR+I0H8ERA2oCCMsCN0
RRRR)Sum<7R=CRs#0kD58IH04E-RI8FMR0Fj
2;S8CMRMoCC0sNCVRH_;IF
VSH_:I4RRHV58IH0>ERR8IH0REq+HRI8A0E2CRoMNCs0RC
RSRRu7)m58IH0+EqI0H8E4A-RI8FMR0Fj<2R=CRs#0kD58IH0+EqI0H8E4A-RI8FMR0Fj
2;SFSVsF_DFIb_:FRVsRRHHIMRHE80qH+I8A0ERR0FI0H8ER-4oCCMsCN0
SSSu7)m5RH2<s=RCD#k0H5I8q0E+8IH0-EA4
2;SMSC8CRoMNCs0VCRFDs_F_FbIS;
CRM8oCCMsCN0R_HVI
4;CRM8NEsO4
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$vR1zRpaHR#
RoRRCsMCH
O5SRRRR8IH0RER:MRH0CCos=R:R;.c
RSRRIRNHE80RH:RMo0CC:sR=.R4;R
SRLRRI0H8ERR:HCM0oRCs:4=R.S
SS
2;RRRRb0Fs5R
SqH:RM0R#8F_Do_HOP0COFNs5I0H8E4R-RI8FMR0Fj
2;RRRRRRRRRRA:H#MR0D8_FOoH_OPC05FsL8IH0-ER4FR8IFM0R;j2
RRRRRRRR)Rum:7RR0FkR8#0_oDFHPO_CFO0sH5I8R0E-84RF0IMF2Rj
RSS2C;
M18Rvazp;N

sHOE00COkRsCODCD_PDCCFDRVvR1zRpaH
#
SMVkOF0HMNROD8IH0REL5MOF#M0N0NRI,LRIRH:RMo0CCRs2skC0sHMRMo0CCHsR#S
SPHNsNCLDRMsO0RR:HCM0o;Cs
CSLo
HMSVSHRL5IRR<=IRN20MEC
SSSs0OMRR:=I;LR
CSSDR#C
SSSs0OMRR:=I;NR
CSSMH8RVS;
S0sCkRsMs0OM;C
SMO8RNHDI8L0E;S

VOkM0MHFRDONI0H8E5NRO#FM00NMR,INRRIL:MRH0CCoss2RCs0kMMRH0CCos#RH
PSSNNsHLRDCs0OMRH:RMo0CC
s;SoLCHSM
SRHV5RIL<I=RN02RE
CMSsSSORM0:I=RN
R;SDSC#
CRSsSSORM0:I=RL
R;SMSC8VRH;S
SskC0ssMRO;M0
MSC8NROD8IH0;EN
O
SF0M#NRM0I0H8E:NRR0HMCsoCRR:=OINDHE80NI5NHE80,IRLHE802S;
O#FM00NMR8IH0REL:MRH0CCos=R:RDONI0H8ENL5I0H8EL,RI0H8E
2;
FSOlMbFCRM0#DlNDDvk0S
SoCCMs5HO
SSSN8IH0:ERR0HMCsoCRS;
SISLHE80RH:RMo0CC;sR
SSSI0H8E:RRR0HMCsoC
2SS;S
Sb0FsRS5
SRSqR:RRRRHMR8#0_oDFHPO_CFO0sI5NHE80-84RF0IMF2Rj;S
SSRARRRR:HRMR#_08DHFoOC_POs0F5HLI8-0E4FR8IFM0R;j2
SSSu7)mRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S
S2S;
CRM8ObFlFMMC0
;
So#HMRNDNk_NG:RRR8#0_oDFHPO_CFO0sH5I8N0E-84RF0IMF2Rj;
RRSo#HMRNDLk_NG:RRR8#0_oDFHPO_CFO0sH5I8L0E-84RF0IMF2Rj;SR
#MHoNsDRCD#k0RR:#_08DHFoOC_POs0F58IH0+ENI0H8E4L-RI8FMR0Fj
2;LHCoM-
S-CRp0R'##bIN
wSQ__IN#_kbIRL:H5VRN8IH0>ER=IRLHE802CRoMNCs0SC
SNN_k<GR=;RN
LSS_GNkRR<=LS;
CRM8oCCMsCN0R_QwI#N_kIb_L
;
S_QwI#L_kIb_NH:RVLR5I0H8ERR>N8IH0RE2oCCMsCN0
NSS_GNkRR<=LS;
SNL_k<GR=;RN
MSC8CRoMNCs0QCRwL_I_b#k_;IN
H
SV4_I:VRHRH5I8L0ER4=R2CRoMNCs0SC
So#HMRNDObFlDCClMR0,0OIFFRlb:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
SLHCoMS
SV_FsDbFF:FRVsRRHHjMRRR0FI0H8E4N-RMoCC0sNCS
SSlOFblDCC5M0H<2R=FRM0_RNN5kGHR2;
CSSMo8RCsMCNR0CV_FsDbFF;S
SSlOFblDCC5M0I0H8E2-4RR<=MRF0Nk_NGH5I8N0E-;42
SSS0OIFFRlb<O=RFDlbCMlC0RR+';4'
sSSCD#k0=R<RhBmea_17m_pt_QBea Bmj)5,HRI8N0E+8IH02ELRCIEMLR5_GNk5Rj2=jR''S2
SCSSDR#C0OIFF;lb

SSS)Sum<7R=CRs#0kD58IH04E-RI8FMR0Fj
2;S8CMRMoCC0sNCVRH_;I4
H
SVj_I:VRHRH5I8L0ER.=R2CRoMNCs0SC
So#HMRNDObFlDCClMR0,0OIFFRlb:0R#8F_Do_HOP0COFIs5HE80NR-48MFI0jFR2S;
LHCoMS
SV_FsDbFF:FRVsRRHHjMRRR0FI0H8E4N-RMoCC0sNCS
SSlOFblDCC5M0H<2R=FRM0_RNN5kGHR2;
CSSMo8RCsMCNR0CV_FsDbFF;S
S0OIFFRlb<O=RFDlbCMlC0RR+';4'
S
SskC#D<0R=mRBh1e_ap7_mBtQ_Be a5m)jN,RI0H8EI+LHE802ERIC5MRLk_NG25jR'=RjN'RML8R_GNk5R42=jR''S2
SCSSDR#C0OIFF5lbI0H8E4N-2RR&0OIFF5lbI0H8E4N-2RR&0OIFFRlbIMECR_5LN5kG4=2RR''4R8NMRNL_kjG52RR='24'
SSSS#CDCIR0FlOFbH5I8N0E-R42&IR0FlOFbRR&'Rj'IMECR_5LN5kG4=2RR''4R8NMRNL_kjG52RR='2j'
SSSS#CDC_RNN5kGI0H8E4N-2RR&Nk_NGH5I8N0E-R42&_RNNRkG;S

Smu)7=R<R#sCk5D0I0H8ER-48MFI0jFR2S;
CRM8oCCMsCN0R_HVI
j;
VSH_:IdRRHV58IH0REL>2R.RMoCC0sNCS
Sl0kD4R:R#DlNDpvzaS
SSCSoMHCsONRlb
R5SSSSSNSSI0H8E>R=R8IH0,EN
SSSSSSSL8IH0=ER>HRI8L0E,S
SSSSSS8IH0RER=I>RHE80
SSSSS2
SbSSFRs0lRNb5S
SSSSSS=qR>_RNN,kG
SSSSSSSA>R=RNL_k
G,SSSSSuSS)Rm7=u>R)
m7SSSS2S;
CRM8oCCMsCN0R_HVI
d;
8CMRDOCDC_DP;CD
