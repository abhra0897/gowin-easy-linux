@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnj-.jRn3qRDDsEHo0s#RCs#CP3C8

RRRNRbsCNl0RCsNC##sM0_NRlC=qR"1)1 a _he_ )zhhim_Whqh1YB
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
R`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MCRCR`MV8H
H
`VV8CRpme_1q1 _)am
h
RDRNI#N$R5@@00C#_bCGsL2RCMoH
RRRRRHV5e`mp _)1_ a1hQtq!pR='R4LRj2LHCoM`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR

Rqq_1)1 a1_qY_hBh  e)h_ziWhmh:_uRR
RNC##s50R!H5f#	kMMMFI5#0C0G_Cb2s22DRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
C
`MV8HRm//eXp_BB] iw_mwR

RCRRMR8
R8CM
C
`MV8HRR//m_epq 11)ma_h



