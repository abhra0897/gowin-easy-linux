@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ha_ )e _izhhhmW"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
`RRHCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0MRC
RM`C8
HV
V`H8RCVm_epq 11)ma_h`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
RRsRbFsbC0q$R1)1 a _he_ )zhhim_WhuR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RJRRkHNDVsHCR>|-Rf!5HM#k	IMFMC50#C0_G2bs2R;
RCRRMs8bFsbC0`$
CHM8V/R/Rpme_]XB _Bim
ww
oRRCsMCN
0C
RRRR#ONCbR5sCFbs_0$0C$b2R
RRRRR`pme_1q1 R)a:CRLoRHM:PRFD#_N#0Cs
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
RRRRRRRRqq_1)1 a _he_ )zhhim_WhuN:R#s#C0sRbFsbC05$Rq 11)ha_ )e _izhhhmW_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
M`C8RHV/m/ReXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lC
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRRRRRRRRv1_q1a )_eh  z)_hmihWuh_:#RN#CklRFbsb0Cs$qR51)1 a _he_ )zhhim_Whu
2;`8CMH/VR/eRmpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
R
RRVRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRRRH5VRm_epB me)q_A1_QBmRh2LHCoMRR:F_PDOCFPsN_L#
HO
RRRRORRFsPC_NJkDHHVC
s:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRJDkNHCVHs22R
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs0J5"kHNDVsHCRPOFC8sC"
2;RRRRR8CMRL//NO#HRPOFCosNCR

RRRRH5VRm_epB me)q_1hYQa_2mhRoLCH:MRRDFP_POFC#s_N0MH$R

RRRRRPOFC0s_C_#0CsGb_NOEM:oC
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjRR&&JDkNHCVHs&R&
RRRRRRRRRRRRRRRRRRRRfR!#L0ND0C5C_#0CsGb2RR22R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsE_ONCMoRPOFC8sC"
2;RRRRR8CMR#//N0MH$FROPNCsoRC
RCRRM
8
CoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
