-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRR:wRRH8GC-HbFMb0RNNO	o5CRQ0M#NHM0N80CRObN	CNoRO8CDNNs0MHF2-
-RRRRRRRRRRRRR-:
-RRRpsHLNRs$RRR:RHaE#NRbOo	NCER#NRDDLOCRFHlbDRC8HFM0RDNRHNLss-$
-RRRRRRRRRRRRRR:Rl#$LHFDODND$NRMlRC8Q   3-
-RRRRRRRRRRRRR-:
-RRR7CCPDCFbsR#:ROqOCCDDseNR]-7paNBRMQ8R R  u(4jnFRWsM	HosRtF
kb-R-RRRRRRRRRR:RR
R--RkRus#bFCRRR:aRRERH#b	NON#oCRV8CH#MCR#LNHLORHsMN$HRVGRC8bMFH0-
-RRRRRRRRRRRRRR:RN0sHE0lCHVORk0MOH#FM
R--RRRRRRRRRRRR:-
-RhRRFR0CRRRRRR:Ra#EHRObN	CNoR$lNRRLClHF8V8HCRR0FHDMOkR8CNH880MHFN8DRN
0N-R-RRRRRRRRRR:RRRCRsJskHCL8R$FR0F,D#R0LkRRH0l0k#RRHMMIFRNO$REoNMCER0C-
-RRRRRRRRRRRRRR:RCCG0sDMNR0HMCNsVORC#F#sRHDlkNF0HMCRLEHNPFFsRVER0C-
-RRRRRRRRRRRRRR:R8OC#s0HbH3FMRRQ0Hb#RCHsl#L#HD0CRF8RN8FROlMlC0N#RMF8/s-
-RRRRRRRRRRRRRR:RNs00H0LkC0#RFER0CNRbOo	NCCR8OsDNNF0HMR#,LRk0MRF00OFREoNMC-
-RRRRRRRRRRRRRR:RF8sRC0DCCMRN$sRFHMoHNDDRH#MCRRFV0RECb	NONRoC8DCON0sNH3FM
R--RRRRRRRRRRRR:aRREbCRNNO	oLCRFR8$lRN$LOCREoNMCF8RMRD$HNMROsOF8ONMCHRI0-E
-RRRRRRRRRRRRRR:RC0ERs0ClF#RVDRBNCk#RR4nF0VRERH##M0N88Ns3-
-RRRRRRRRRRRRR-:
--R--------------------------------------------------------------------
-)RfC#PHH:FMR.4.j
Rf-f-R7CN0:jR.jjU-cj-4R:4(4jn:gjR+gRdj5kaE,jR4RsqbRj.jUf2R
R----------------------------------------------------------------------
H
DLssN$ RQ R ;RR--oCCMs#HORDLCFsIRCsNsNCMo8FRVsCR#OHks0s$RCFN#M
#
b	NONRoCVCHG8	_bo#RHRIMCR Q  H3VG_C8oCCMs_HOb
	oRCRoMHCsONRlb
R5RRRRVCHG8P_FCDsVF#I_0C$DRR=>Q   3GVHCV8_D0FN_b0$CV#3H8GC_0#Nk0sNCR,
RVRRH8GC_NoksL8_HR0#RRRR=d>R,R
RRHRVG_C8sMFk80_#$RDCR=RR> RQ V 3H8GC_FVDN00_$#bC3GVHCs8_F8kM,R
RRFRM_sINMoHMRRRRRRRRR=RR>NRVD
#CRRRR2
;

