--$Header: //synplicity/mapgw/designware/dw06.vhd#1 $
@E---------------------------------------------------------------------------------------------------

---w-RHRDCRRRRR:RRRj8InE3P8-
-R#7CHRoMRRRRRB:RFNM0HRM#4LURNO#HR#7CHWoMNRsCObFlFMMC0
#R-B-RFNlbMR$RR:RRRM1$bODHHR0$Q3MO
R--7CN0RRRRRRRR:kRqo6R.,jR.j-U
-kRq0sEFRRRRRRR:1PCDN)lR
R--e#CsHRFMRRRR:3Rd4-
-
---------------------------------------------------------------------------------------------------
H
DLssN$ RQ 8 ,I;jdR#
kCIR8j8d3I_jdObFlFMMC0N#3D
D;kR#CQ   38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;#
kCCRHC#C30D8_FOoH_HNs0NE3D
D;
M
C0$H0R_7WNl#$VFHV__#48HVR#S
SoCCMsRHO5S
SS08NNM_H_8IH0:ESRaQh )t RR:=US;
SNS80FN_kI0_HE80SQ:Rhta  :)R=nR4;S
SSb8C0SERSRS:Q hatR ):U=R;RSR
SSSC_sslCF8R:SSRaQh )t RR:=4S;
S#Ss0F_l8SCS:hRQa  t)=R:R
4;SLSS$_0CFCs8s:SSRaQh )t RR:=jS
SS
2;SFSbs50R
RSSRORRDR	RRSSS:MRHR0R#8F_Do;HO
SSSs_#0MSRRSRS:HRMR#_08DHFoOS;
SkSb#sE_CMJ_R:RSRRHMR8#0_oDFH
O;SVSSDEk#_SMSSH:RM#RR0D8_FOoH;S
SSbbF_JsC_RMRRRS:HRMR#_08DHFoOS;
SHS8NMo_RSRS:MRHR0R#8F_Do;HO
SSS8NN0_RHMSRS:HRMR#_08DHFoOC_POs0F508NNM_H_8IH04E-RI8FMR0Fj
2;SNSSCC_DPRCDRRRRR:RRRRHMR8#0_oDFHPO_CFO0s55RR0LH_8IH08E5CEb02RR-482RF0IMFRRj2S;
SVSN_s0ECS#ESH:RM#RR0D8_FOoH_OPC05FsRL5RHI0_HE805b8C0RE2-2R4RI8FMR0Fj;R2SS
SSbCl0R$RS:SSR0FkR8#0_oDFH
O;SNSSD#lF0l_CbS0$:kRF00R#8F_Do;HO
SSSEVND_DVkDSRS:kRF00R#8F_Do;HO
SSSNFDl#V0_kRDDSF:Rk#0R0D8_FOoH;S
SSDVkDSRRSRS:FRk0#_08DHFoOS;
SNSslk_VDSDS:kRF00R#8F_Do;HO
SSSCFsssSRRSRS:FRk0#_08DHFoOS;
SNSbsI0_8SSS:kRF00R#8F_Do;HO
SSS8NN0_0FkSRS:FRk0#_08DHFoOC_POs0F508NNk_F0H_I8-0E4FR8IFM0RSj2
SSSSS
SS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_$N#lVVHF4_#_R8V:MRC0$H0RRH#"NIC	
";
MSC8WR7_$N#lVVHF4_#_;8V
NR
sHOE00COkRsC#k0sOF0RVWR7_$N#lVVHF4_#_R8VH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0R#s0kORN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRs#0kRO0:sRNO0EHCkO0sHCR#sR0k
C;SLR
CMoH
M
C80R#s0kO;



----------------------------------------------------------------------------D-
HNLssQ$R ,  8dIj;kR
#8CRI3jd8dIj_lOFbCFMM30#N;DD
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_#kMHCoM8D3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
M
C0$H0R_7WNl#$VFHV__#4#HVR#S
SoCCMsRHO5S
SS08NNM_H_8IH0:ESRaQh )t RR:=.
c;S8SSN_0NF_k0I0H8ERS:Q hatR ):U=R;S
SSb8C0SERSRS:Q hatR ):U=R;RSR
SSSNDC_CDPCRRRRSQ:Rhta  :)R=;Rc
SSSNDV_CDPCRSRRRRRR:hRQa  t)=R:R
c;SCSSsls_FR8CSRS:Q hatR ):4=R;S
SS0s#_8lFC:SSRaQh )t RR:=4S;
S$SL0FC_ss8CSRS:Q hatR ):j=R
SSS2S;
SsbF0
R5SbSSk_#Es_CJMSRR:MRHR0R#8F_Do;HO
SSSb_Fbs_CJMRRRSH:RM#RR0D8_FOoH;
SRS8SSN_0NHSMRSH:RM#RR0D8_FOoH_OPC05Fs8NN0__HMI0H8ER-48MFI0jFR2S;
SDSVk_#EMSSS:MRHR0R#8F_Do;HO
SSS8NN0_0FkSRS:FRk0#_08DHFoOC_POs0F508NNk_F0H_I8-0E4FR8IFM0R;j2SS
SSlsN_DVkD:SSR0FkR8#0_oDFH
O;SbSSN_s0IS8SSF:Rk#0R0D8_FOoH;S
SSN8HoR_MR:SSRRHMR8#0_oDFH
O;SOSSDR	RRSSS:MRHR0R#8F_Do;HO
SSSs_#0MSRRSRS:HRMR#_08DHFoOS;
SkSVDRDRS:SSR0FkR8#0_oDFH
O;SNSSD#lF0k_VDSDR:kRF00R#8F_Do;HO
SSSEVND_DVkDSRS:kRF00R#8F_Do;HO
SSSNFDl#C0_l$b0SF:Rk#0R0D8_FOoH;S
SSbCl0R$RS:SSR0FkR8#0_oDFH
O;SCSSsssFRSRSSF:Rk#0R0D8_FOoH
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7WNl#$VFHV__#4#:VRR0CMHR0$H"#RI	CN"
;
S8CMR_8INl#$VFHV__#4#
V;Rs
NO0EHCkO0s#CR0Osk0VRFR_7WNl#$VFHV__#4#HVR#-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRs#0kRO0:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFV#k0sO:0RRONsECH0Os0kC#RHRk0sCS;

oLCH
MR
M
C80R#s0kO;S


-
--------------------------------------------------------------------------
--DsHLNRs$Q   ,j8Id
;R-#-kCIR8j8n3I_jnObFlFMMC0N#3D
D;kR#C8dIj3j8IdF_OlMbFC#M03DND;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;


CHM007$RWH_VV#F_4V_#R
H#oCCMsRHO5S
SS8IH0SERRQ:Rhta  :)R=;RU
SSS80CbERRS:hRQa  t)=R:R
c;SNSSCC_DPRCD:hRQa  t)=R:R
4;SNSSVC_DPRCD:hRQa  t)=R:R
4;SCSSsls_FR8C:hRQa  t)=R:R
j;SsSS#l0_FR8C:hRQa  t)=R:RSj
RSRRS
2;b0FsRb5
k_#Es_CJM:RSRRHM#_08DHFoOb;
Fsb_CMJ_R:RSRRHM#_08DHFoO8;
H_NoM:SSRRHM#_08DHFoOO;
DS	RSH:RM0R#8F_Do;HO
0s#_SMS:MRHR8#0_oDFH
O;8NN0_RHMRRRR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
DVkD:SSR0FkR8#0_oDFH
O;NFDl#V0_kSDD:kRF00R#8F_Do;HO
DENVk_VD:DSR0FkR8#0_oDFH
O;NFDl#C0_l$b0:kRF00R#8F_Do;HO
bCl0S$S:kRF00R#8F_Do;HO
sCsFSsS:kRF00R#8F_Do;HO
08NNk_F0RRRRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_VV#F_4V_#RC:RM00H$#RHRC"IN;	"
8CMR_7WVFHV__#4#
V;
N

sHOE00COkRsCsR0DF7VRWH_VV#F_4V_#R
H#
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;

oLCH
MSSM
C80RsD
;

-
--------------------------------------------------------------------------
--
LDHs$NsR Q  I,8jRd;
Ck#Rj8IdI38jOd_FFlbM0CM#D3NDk;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;

0CMHR0$7VW_H_VF#84_V#RH
MoCCOsHRS5
Sb8C0RERRRR:Q hatR ):U=R;S
SI0H8ERRRRQ:Rhta  :)R=;RcSS
SC_sslCF8RQ:Rhta  :)R=;Rj
sSS#l0_FR8C:hRQa  t)=R:RSj
RSRRS
2;b0FsRO5
DS	RSH:RM0R#8F_Do;HO
0s#_SMS:MRHR8#0_oDFH
O;bEk#_JsC_SMR:MRHR8#0_oDFH
O;b_Fbs_CJMSRR:MRHR8#0_oDFH
O;8oHN_SMS:MRHR8#0_oDFH
O;NDC_CDPCRRRR:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;N0V_E#sCERRR:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;8NN0_RHMRRRR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
bCl0S$S:kRF00R#8F_Do;HO
lNDF_#0C0lb$F:Rk#0R0D8_FOoH;N
EDVV_kSDD:kRF00R#8F_Do;HO
DVkD:SSR0FkR8#0_oDFH
O;NFDl#V0_kSDD:kRF00R#8F_Do;HO
sCsFSsS:kRF00R#8F_Do;HO
08NNk_F0RRRRF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2;
2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWH_VV#F_4V_8RC:RM00H$#RHRC"IN;	"
M
C8WR7_VVHF4_#_;8V



NEsOHO0C0CksRDs0RRFV7VW_H_VF#84_V#RH
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
oLCHSMS
SSS
8CMRDs0;-

------------------------------------------------------------------------------------
H
DLssN$ RQ 8 ,I;jd
Ck#R Q  03#8F_Do_HO4c4n3DND;#
kC RQ # 30D8_FOoH_HNs0NE3D
D;kR#CQ   38#0_oDFHkO_Mo#HM3C8N;DD
Ck#Rj8IdI38jOd_FFlbM0CM#D3ND
;
CHM007$RWH_VV#F_.V_#R
H#oCCMs5HORS
SI0H8ESRS:hRQa  t)=R:R
U;SCS8bR0ESRS:Q hatR ):U=R;S
SbEk#__NCDRPD:hRQa  t)=R:R
.;SkSb#NE_VP_DDRR:Q hatR ):.=R;S
Sb_FbNDC_PRDR:hRQa  t)=R:R
.;SFSbbV_N_DDPRRR:Q hatR ):.=R;S
SC_sslCF8RRS:Q hatR ):j=R;S
SbEk#_M#$O:RSRaQh )t RR:=.S;
SbbF_M#$O:RSRaQh )t RR:=.S;
S0s#_8lFC:RSRaQh )t RR:=dSR
SSS
S;S2SSR
SSS

R
RRRRRRsbF0RR5
RRRRRRRRRRRR	OD_#bkERRS:MRHR8#0_oDFH;OR
SSSO_D	bSFbRRRRRH:RM0R#8F_Do;HO
RRRRRRRR#Ss0R_MSRRS:MRHR8#0_oDFH;OR
RRRRRRRRkSb#sE_CMJ_SRR:H#MR0D8_FOoHRS;
SFSbbC_sJS_MRH:RM0R#8F_DoRHO;S
SS08NNM_HS:SRRRHM#_08DHFoOC_POs0FR55RI0H8ERR-482RF0IMFRRj2S;
SkSb#CE_l$b0SRR:FRk0#_08DHFoOS;
SkSb#NE_C:SRR0FkR8#0_oDFH
O;SbSSk_#EERVS:kRF00R#8F_Do;HO
SSSbEk#_SNVRF:Rk#0R0D8_FOoH;S
SS#bkEk_VDRDS:kRF00R#8F_Do;HO
SSSbEk#_sCsFRsS:kRF00R#8F_Do;HO
SSSb_FbC0lb$:SRR0FkR8#0_oDFH
O;SbSSFNb_C:SRR0FkR8#0_oDFH
O;SbSSFEb_V:SRR0FkR8#0_oDFH
O;SbSSFNb_V:SRR0FkR8#0_oDFH
O;SbSSFVb_kSDDRF:Rk#0R0D8_FOoH;R
SSFSbbs_CsSFsRF:Rk#0R0D8_FOoH;S
SS08NNk_F0RRRRRR:FRk0#_08DHFoOC_POs0FRI55HE80R4-RR82RF0IMFRRj2S

S
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_VVHF._#_R#V:MRC0$H0RRH#"NIC	
";SM
C8IR8_VVHF._#_;#V
s
NO0EHCkO0s#CR0Osk0VRFR_8IVFHV__#.#HVR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0R#s0kORN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRs#0kRO0:sRNO0EHCkO0sHCR#sR0k
C;


SLHCoM
RR
8CMRs#0k;O0



-=-=====================================CHM00N$RMN8RsHOE00COkRsCVRFs8#I_0	NO=============================D

HNLssH$RC,CC8nIj,j8Idk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#8CRI3jn8nIj_lOFbCFMM30#N;DD
Ck#Rj8IdI38jOd_FFlbM0CM#D3ND
;

SS
CHM007$RW0_#NRO	HS#
SMoCCOsHRS5
SHSI8R0ESRR:Q hatR ):U=R;S
SSb8C0SERRQ:Rhta  :)R=;RU
SSSC_sslCF8RQ:Rhta  :)R=;Rj
SSSs_#0lCF8RQ:Rhta  :)R=
RjS2SS;S
Sb0FsRS5
SDSO	SRS:MRHR8#0_oDFH
O;SsSS#M0_R:SSRRHM#_08DHFoOS;
SkSb#sE_CMJ_RRR:H#MR0D8_FOoH;S
SSbbF_JsC_SMR:MRHR8#0_oDFH
O;S8SSN_0NHSMR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
SSSC0lb$SRS:kRF00R#8F_Do;HO
SSSVDkDR:SSR0FkR8#0_oDFH
O;SCSSsssFR:SSR0FkR8#0_oDFH
O;S8SSN_0NFRk0SF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S
SS
2;
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_N#0O:	RR0CMHR0$H"#RI	CN"
;
S8CMR_7W#O0N	
R;
N
SsHOE00COkRsCsR0DF7VRW0_#NRO	H
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;

SSC
Lo
HM
M
C80RsD
;

=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFR_7W)_qv)qW__w7wR========================
=

LDHs$NsR Q  I,8jRn;
Ck#R Q  03#8F_po_HO4c4n3DqD;kR
#QCR 3  #_08pHFoOM_k#MHoCq83DRD;R#
kCIR8j8n3I_jnObFlFMMC0N#3D
D;
0CMHR0$7sW_Nsl_I__N8RVVHS#
SMoCCOsHRS5
SNS80IN_HE80RQ:Rhta  :)R=;RU
SSS80CbERRRR:RRRaQh )t RR:=US;
S#Ss0F_l8RCRRQ:Rhta  :)R=
RjS2SS;S
Sb0FsRS5
S#Ss0R_MRRRRR:RRRRHMR8#0_oDFH
O;SOSS#R_MRRRRRRRR:MRHR0R#8F_Do;HO
SSSIMs_RRRRRRRRRH:RM#RR0D8_FOoH;
SRS0SSC_#0lCF8RRRR:MRHR0R#8F_Do;HO
SSS00C#_	ODRRRRRH:RM#RR0D8_FOoH;S
SS_sINs88RRRRRRR:HRMR#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SNS80HN_MRRRR:RRRRHMR8#0_oDFHPO_CFO0sN580IN_HE80-84RF0IMF2Rj;S
SS08NNk_F0RRRRRR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0RSj2
SSS2
;
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7Ws_NlsNI__V8VRC:RM00H$#RHRC"IN;	"
M
C8WR7_lsN__sINV_8VR;RR


NEsOHO0C0CksRDs0RRFV7sW_Nsl_I__N8RVVH
#
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;

=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFR_7W)_qv)qW__apq=========================D

HNLssQ$R ,  8nIj;kR
#QCR 3  #_08pHFoO4_4nqc3DRD;
Ck#R Q  03#8F_po_HOkHM#o8MC3DqD;
RRkR#C8nIj3j8InF_OlMbFC#M03DND;


CHM007$RWN_slI_s_DN_NH0R#S
SoCCMsRHO5S
SS08NNH_I8R0E:hRQa  t)=R:R
g;S8SSCEb0RRRRRRR:Q hatR ):4=RcS;
S#Ss0F_l8RCRRQ:Rhta  :)R=
RjS2SS;S
Sb0FsRS5
S#Ss0R_MSRRR:MRHR0R#8F_Do;HO
SSSOM#_RRSRRH:RM#RR0D8_FOoH;S
SS_IsMRRRRRRR:MRHR0R#8F_Do;HO
SSSsNI_8R8sR:RRRRHMR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;S8SSN_0NHRMRRRR:HRMR#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R;j2
SSS8NN0_0FkR:RRR0FkR8#0_oDFHPO_CFO0sN580IN_HE80-84RF0IMF2Rj
SSS2-;
-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7sW_Nsl_I__NDRN0:MRC0$H0RRH#"NIC	
";
8CMR_7Ws_NlsNI__0DNRS;R
s
NO0EHCkO0ssCR0FDRVWR7_lsN__sINN_D0HRR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
M
C80RsD
;

-R-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7_v)q_W)__7q_w=w======================
==
H
DLssN$ RQ 8 ,I;jnR#
kC RQ 1 30p8_FOoH_n44cD3qD
;RkR#CQ   3810_opFHkO_Mo1HM3C8q;DDRkR
#8CRI3jn8nIj_lOFbCFMM30#N;DD
M
C0$H0R_7Ws_Nls__INV_8V#RH
oSSCsMCH5OR
SSS8NN0_8IH0:ERRaQh )t RR:=cS;
SCS8bR0ERRRRRQ:Rhta  :)R=;RU
SSSs_#0lCF8R:RRRaQh )t RR:=jS
SSS2;SS
Sb0FsRS5
S#Ss0R_MRRRRRH:RM#RR0D8_FOoH;S
SS_O#MRRRRRRR:MRHR0R#8F_Do;HO
SSSIMs_RRRRR:RRRRHMR8#0_oDFH
O;S0SSC_#0lCF8RRR:HRMR#_08DHFoOS;
SCS0#O0_DR	RRH:RM#RR0D8_FOoH;S
SS_s8Ns88RRRR:MRHR0R#8F_Do_HOP0COFLs5HI0_HE80RC58b20E-84RF0IMF2Rj;S
SS_IsNs88RRRR:MRHR0R#8F_Do_HOP0COFLs5HI0_HE80RC58b20E-84RF0IMF2Rj;S
SS08NNM_HRRRR:MRHR0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2S;
SNS80FN_kR0RRF:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0Fj
2RS2SS;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWN_sl__sI__N8RVV:MRC0$H0RRH#"NIC	
";
8CMR_7Ws_Nls__INV_8VRR;
s
NO0EHCkO0ssCR0FDRVWR7_lsN_Is__8N_VRVRH
#R
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIs
CRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoN;
0H0sLCk0RM#$_HLkDM0H_R8kFsVR0:DRRONsECH0Os0kC#RHRC"IN;	"
-R
-FRwsHR#MCoDRk#FsROC7RW,NEsOHO0C0CksRF#EkRD8L8CRk$ll
0N0skHL0#CR$LM_D	NO_GLFRL:RFCFDN
M;Ns00H0LkC$R#MD_LN_O	LRFGFsVR0:DRRONsECH0Os0kC#RHRk0sC
;
LHCoM

RCRM8s;0D



-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs7)W_q)v__qW__apq=========================D

HNLssQ$R ,  8nIj;kR
#QCR 3  #_08pHFoO4_4nqc3DRD;
Ck#R Q  03#8F_po_HOkHM#o8MC3DqD;kR
#8CRI3jn8nIj_lOFbCFMM30#N;DD
C

M00H$WR7_lsN_Is__DN_NH0R#C
oMHCsO
R58NN0_8IH0:ERRaQh )t RR:=U8;
CEb0RQ:Rhta  :)R=nR4;#
s0F_l8:CRRaQh )t RR:=j;
2
F
bs50R
0s#_:MRRRHM#_08DHFoOO;
#R_M:MRHR8#0_oDFH
O;IMs_RH:RM0R#8F_Do;HO
_s8Ns88RH:RM0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
_IsNs88RH:RM0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
08NNM_HRH:RM0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR28;
N_0NFRk0:kRF00R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2;
2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_lsN_Is__DN_N:0RR0CMHR0$H"#RI	CN"
;
CRM87sW_Nsl__NI__0DNR
;R
ONsECH0Os0kC0RsDVRFR_7Ws_Nls__INN_D0#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
C
Lo
HM
8CMRDs0;S
SS
S

-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7_v)q__.)W__q7=ww========================
D

HNLssQ$R ,  8nIj;kR
#QCR 3  1_08pHFoO4_4nqc3DRD;
Ck#R Q  0318F_po_HOkHM#o8MC3DqD;
RRkR#C8nIj3j8InF_OlMbFC#M03DND;C

M00H$WR7_lsN__.sI__N8RVVHS#SSRSSRSR
SMoCCOsHRS5
SNS80IN_HE80RQ:Rhta  :)R=;Rc
SSS80CbERRRR:RRRaQh )t RR:=cS;
S#Ss0F_l8RCRRQ:Rhta  :)R=
RjS2SS;SS
SsbF0
R5SsSS#M0_RRRRRRRR:MRHR0R#8F_Do;HO
SSSOM#_RRRRRRRRRH:RM#RR0D8_FOoH;S
SS_IsMRRRRRRRRRR:HRMR#_08DHFoOS;
SCS0#l0_FR8CR:RRRRHMR8#0_oDFH
O;S0SSC_#0ORD	RRRR:MRHR0R#8F_Do;HO
SSSs_84Ns88RRRRRH:RM#RR0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS.s8_8N8sRRRRRR:HRMR#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SsSI_8N8sRRRR:RRRRHMR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;S8SSN_0NHRMRRRRR:MRHR0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2S;
SNS80sN_8F4_k:0RR0FkR8#0_oDFHPO_CFO0sN580IN_HE80-84RF0IMF2Rj;S
SS08NN8_s.k_F0RR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R
j2S2SS;-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNs
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;RRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8RRFV7sW_N.l_s__INV_8VRR:CHM00H$R#IR"C"N	;C

M78RWN_sls_._NI__V8VRR;RS
S
NEsOHO0C0CksRDs0RRFV7sW_N.l_s__INV_8VHRR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;L

CMoH
CR
Ms8R0
D;




-R
-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRWq_)v)_._qW__apq=========================H
DLssN$ RQ 8 ,I;jnR#
kC RQ # 30p8_FOoH_n44cD3qD
;RkR#CQ   38#0_opFHkO_Mo#HM3C8q;DDRkR
#8CRI3jn8nIj_lOFbCFMM30#N;DD
C

M00H$WR7_lsN__.sI__NDRN0HS#
SMoCCOsHRS5
SNS80IN_HE80RQ:Rhta  :)R=.R4;S
SSb8C0RERRRRR:hRQa  t)=R:R;4c
SSSs_#0lCF8R:RRRaQh )t RR:=4S
SS
2;SFSbs50R
SSSs_#0MRRSRRR:HRMR#_08DHFoOS;
S#SO_SMRR:RRRRHMR8#0_oDFH
O;SISSsR_MRRRRRRR:HRMR#_08DHFoOS;
S8Ss48_N8RsRRRR:HRMR#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
S8Ss.8_N8RsRRRR:HRMR#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SsSI_8N8sRRRRH:RM#RR0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS08NNM_HRRRR:MRHR0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2S;
SNS80sN_8F4_kR0RRF:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0Fj
2;S8SSN_0Ns_8.FRk0RRR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R
j2S2SS;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWN_sls_._NI__0DNRC:RM00H$#RHRC"IN;	"
M
C8WR7_lsN__.sI__NDRN0;N

sHOE00COkRsCsR0DF7VRWN_sls_._NI__0DNR#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC
L

CMoH
C

Ms8R0
D;R-S
-========================================C==M00H$MRN8sRNO0EHCkO0sVCRF7sRWq_)vW_)_71_wRwSR========================
=
DsHLNRs$Q   ,j8In
;RkR#CQ   3810_opFH4O_43ncq;DDR#
kC RQ 1 30p8_FOoH_#kMHCoM8D3qDR;R
Ck#Rj8InI38jOn_FFlbM0CM#D3ND
;

0CMHR0$7sW_Nsl_I__#8RVVHS#
SMoCCOsHRS5
SNS80IN_HE80RQ:Rhta  :)R=;Rc
SSS80CbERRSRRR:Q hatR ):c=R;S
SS0s#_8lFCRRR:hRQa  t)=R:RSj
S;S2
bSSFRs05S
SS	ODR:SSRRHM#_08DHFoOS;
S#Ss0R_MSRS:H#MR0D8_FOoH;S
SS_O#MSRS:MRHR8#0_oDFH
O;SISSsR_MSRS:H#MR0D8_FOoH;S
SS_sINs88RRS:H#MR0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS08NNM_HRRS:H#MR0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0Fj
2;S8SSN_0NFRk0SF:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0FjS2
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_lsN__sI#V_8VRR:CHM00H$R#IR"C"N	;C

M78RWN_slI_s_8#_V
V;
ONsECH0Os0kC0RsDVRFR_7Ws_Nls#I__V8VRRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
C
LoRHM
M
C80RsDRR;
-
-=========================================M=C0$H0R8NMRONsECH0Os0kCFRVsWR7_v)q__)W1q_pa=RR========================
H
DLssN$ RQ 8 ,I;jnR#
kC RQ 1 30p8_FOoH_n44cD3qD
;RkR#CQ   3810_opFHkO_Mo1HM3C8q;DDRkR
#8CRI3jn8nIj_lOFbCFMM30#N;DD
M
C0$H0R_7Ws_Nls#I__0DNRRH#
oSSCsMCH5ORRS
SS08NNH_I8R0E:hRQa  t)=R:R
c;S8SSCEb0RRRRRRR:Q hatR ):c=R
RSSR2RR;
SSSFSbsR05
SSSORD	RRRRR:RRRRHMR8#0_oDFH
O;SOSS#R_MRRRRRRR:HRMR#_08DHFoOS;
SsSI_RMRRRRRRH:RM#RR0D8_FOoH;S
SS_sINs88RRRR:MRHR0R#8F_Do_HOP0COF5sRL_H0I0H8E8R5CEb02R-48MFI0jFR2S;
SNS80HN_MRRRRH:RM#RR0D8_FOoH_OPC0RFs508NNH_I8-0E4FR8IFM0R;j2
SSS8NN0_0FkR:RRR0FkR8#0_oDFHPO_CFO0s8R5N_0NI0H8ER-48MFI0jFR2SS
S;S2
R--Ns00H0LkCCR8OsDNNF0HMFRVsHR#MCoDRk#FsROC8HC#oNMIsRC
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;R
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8FkRVWR7_lsN__sI#N_D0RR:CHM00H$R#IR"C"N	;C

M78RWN_slI_s_D#_N;0RRN

sHOE00COkRsCsR0DF8VRIN_slI_s_D#_NH0R#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;

R
oLCH
M

8CMRDs0;



=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFR_7W)_qv)__W1w_7w=RR========================
H
DLssN$ RQ 8 ,I;jnR#
kC RQ 1 30p8_FOoH_n44cD3qD
;RkR#CQ   3810_opFHkO_Mo#HM3C8q;DDRkR
#8CRI3jn8nIj_lOFbCFMM30#N;DDR


CHM007$RWN_sl__sI__#8RVVHS#
SMoCCOsHRS5
SNS80IN_HE80RQ:Rhta  :)R=;RU
SSS80CbERRSRRR:Q hatR ):U=R;S
SS0s#_8lFCRRR:hRQa  t)=R:RSj
S;S2
bSSFRs05S
SS	ODRSSS:MRHR8#0_oDFH
O;SsSS#M0_RSSS:MRHR8#0_oDFH
O;SOSS#R_MS:SSRRHM#_08DHFoOS;
SsSI_SMRSRS:H#MR0D8_FOoH;S
SS_s8Ns88R:SSRRHM#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SsSI_8N8sSRS:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;S8SSN_0NHSMRSH:RM0R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2S;
SNS80FN_kS0R:kRF00R#8F_Do_HOP0COF8s5N_0NI0H8ER-48MFI0jFR2S
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7Ws_Nls__I#V_8VRR:CHM00H$R#IR"C"N	;C
SM78RWN_sl__sI__#8;VV
s
NO0EHCkO0ssCR0FDRVIR8_lsN_Is__8#_VHVR#
R
-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCNR
0H0sLCk0RM#$_HLkDM0H_R8k:0R#soHM;0
N0LsHkR0C#_$MLDkH0_HM8FkRV0RsDRR:NEsOHO0C0CksRRH#"NIC	
";R-
-RswFRM#HoRDC#sFkO7CRWN,RsHOE00COkRsC#kEFDL8RCkR8l
l$Ns00H0LkC$R#MD_LN_O	LRFG:FRLFNDCMN;
0H0sLCk0RM#$_NLDOL	_FFGRV0RsDRR:NEsOHO0C0CksRRH#0Csk;S


oLCH
M
CRM8sR0D;


-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs7)W_q)v__1W__apqR=R======================
==DsHLNRs$Q   ,j8In
;RkR#CQ   3810_opFH4O_43ncq;DDR#
kC RQ 1 30p8_FOoH_#kMHCoM8D3qDR;R
Ck#R Q  0318F_po_HON0sHED3qDR;R
Ck#Rj8InI38jOn_FFlbM0CM#D3ND
;R
M
C0$H0R_7Ws_Nls__I#N_D0#RHRS
SoCCMsRHO5SR
SNS80IN_HE80RQ:Rhta  :)R=;Rc
SSS80CbERRRR:RRRaQh )t RR:=US
SSS2;SS
Sb0FsR
5RSsSS88_N8RsR:MRHR0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
SSSINs_8R8sRH:RM#RR0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS08NNM_HRRR:HRMR#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R;j2
SSSOSD	SRR:HRMR#_08DHFoOS;
S#SO_RMRR:RRRRHMR8#0_oDFH
O;SISSsS_MRH:RM#RR0D8_FOoH;S
SS08NNk_F0RR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R
j2S2SS;-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWN_sl__sI__#DRN0:MRC0$H0RRH#"NIC	
";CRM87sW_Nsl__#I__0DNR
;R
ONsECH0Os0kC0RsDVRFR_7Ws_Nls__I#N_D0#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC

S
LHCoM
R
CRM8s;0D




=--=========================================0CMHR0$NRM8NEsOHO0C0CksRsVFR_7W)_qv.W)__71_wRwR=========================D

HNLssQ$R ,  8nIj;kR
#QCR 3  1_08pHFoO4_4nqc3DRD;
Ck#R Q  0318F_po_HOkHM#o8MC3DqD;
RRkR#C8nIj3j8InF_OlMbFC#M03DND;
R

0CMHR0$7sW_N.l_s__I#V_8V#RH
oSSCsMCH5OR
SSS8NN0_8IH0:ERRaQh )t RR:=US;
SCS8bR0ESRRR:hRQa  t)=R:R
U;SsSS#l0_FR8CRRR:Q hatR ):j=R
SSS2S;
SsbF0
R5SOSSDS	RSRS:H#MR0D8_FOoH;S
SS0s#_SMRSRS:H#MR0D8_FOoH;S
SS_O#MSRSSH:RM0R#8F_Do;HO
SSSIMs_RSSS:MRHR8#0_oDFH
O;SsSS8N4_8R8sSRS:H#MR0D8_FOoH_OPC05FsL_H0I0H8EC58b20E-84RF0IMF2Rj;S
SS.s8_8N8sSRS:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;SISSs8_N8SsRSH:RM0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
SSS8NN0_RHMSRS:H#MR0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0Fj
2;S8SSN_0Ns_84FRk0SF:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0Fj
2;S8SSN_0Ns_8.FRk0SF:Rk#0R0D8_FOoH_OPC05Fs8NN0_8IH04E-RI8FMR0FjS2
S;S2
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMN
sCRRRRRRRRNs00H0LkC$R#Mk_LHHD0Mk_8R#:R0MsHoR;
RRRRRNRR0H0sLCk0RM#$_HLkDM0H_R8kF7VRWN_sls_._#I__V8VRC:RM00H$#RHRC"IN;	"
C
SM78RWN_sls_._#I__V8V;N

sHOE00COkRsCsR0DF8VRIN_sls_._#I__V8VRRH#
-
-R0N0skHL08CRCNODsHN0FVMRF#sRHDMoCFR#kCsOR#8CHIoMNRsC
0N0skHL0#CR$LM_k0HDH8M_kRR:#H0sM
o;Ns00H0LkC$R#Mk_LHHD0Mk_8RRFVsR0D:sRNO0EHCkO0sHCR#IR"C"N	;

R-w-RF#sRHDMoCFR#kCsOR,7WRONsECH0Os0kCER#F8kDRRLC8lkl$0
N0LsHkR0C#_$MLODN	F_LGRR:LDFFC;NM
0N0skHL0#CR$LM_D	NO_GLFRRFVsR0D:sRNO0EHCkO0sHCR#sR0k
C;
LS
CMoHR

SSM
C80RsD
R;



-=-=========================================CHM00N$RMN8RsHOE00COkRsCVRFs7)W_q.v_)__W1q_pa========================D=
HNLssQ$R ,  8nIj;kR
#QCR 3  1_08pHFoO4_4nqc3DRD;
Ck#R Q  0318F_po_HOkHM#o8MC3DqD;
RRkR#CQ   3810_opFHNO_sEH03DqD;kR
#8CRI3jn8nIj_lOFbCFMM30#N;DDRC

M00H$WR7_lsN__.sI__#DRN0HS#
SMoCCOsHR
5RS8SSN_0NI0H8ERR:Q hatR ):U=R;S
SSb8C0RERRRRR:hRQa  t)=R:RSU
S;S2S
SSSFSbs50RRS
SS	ODRRSSRH:RM0R#8F_Do;HO
SSSOM#_RRRRS:RRRRHM#_08DHFoOS;
SsSI_RMRRRRSRH:RM0R#8F_Do;HO
SSSs_84Ns88RRSR:MRHR8#0_oDFHPO_CFO0sH5L0H_I850E80CbE42-RI8FMR0Fj
2;SsSS8N._8R8sS:RRRRHM#_08DHFoOC_POs0F50LH_8IH08E5CEb02R-48MFI0jFR2S;
SsSI_8N8sRSSRH:RM0R#8F_Do_HOP0COFLs5HI0_HE805b8C0-E24FR8IFM0R;j2
SSS8NN0_RHMS:RRRRHM#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R;j2
SSS8NN0_4s8_0FkRRR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0R;j2
SSS8NN0_.s8_0FkRRR:FRk0#_08DHFoOC_POs0F508NNH_I8-0E4FR8IFM0RRj2RRSRRS
SS
2;-N-R0H0sLCk0RO8CDNNs0MHFRsVFRM#HoRDC#sFkO8CRCo#HMsINCR
RRRRRR0RN0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
RRRRRRRR0N0skHL0#CR$LM_k0HDH8M_kVRFR_7Ws_Nl.Is__D#_N:0RR0CMHR0$H"#RI	CN"
;
CRM87sW_N.l_s__I#N_D0
;
NEsOHO0C0CksRDs0RRFV7sW_N.l_s__I#N_D0#RHR-

-0RN0LsHkR0C8DCON0sNHRFMVRFs#oHMD#CRFOksCCR8#MHoICNsR0
N0LsHkR0C#_$MLDkH0_HM8:kRRs#0H;Mo
0N0skHL0#CR$LM_k0HDH8M_kVRFRDs0RN:RsHOE00COkRsCH"#RI	CN"R;

R--wRFs#oHMD#CRFOksCWR7,sRNO0EHCkO0s#CREDFk8CRLRl8klN$
0H0sLCk0RM#$_NLDOL	_F:GRRFLFDMCN;0
N0LsHkR0C#_$MLODN	F_LGVRFRDs0RN:RsHOE00COkRsCH0#Rs;kC


SLHCoMSR

CS
Ms8R0RD;




