--=============================== entity and architecture dw_div===============================
@E-

-------------------------------------------------------------------------------------------------
-----
-HRa0RDCRRRRRRR:78W_H-P
-CR7#MHoRRRRRRR:78W_H-P
-kRq0sEFRRRRRRR:1PCDN)lRR]/RN#sHERRvi-
-RlBFb$NMRRRRR1:R$DMbH0OH$FR1VN0IsQCRMN8HR0uP30Rp8-3
--
---------------------------------------------------------------------------------------------------
-R#7CObsH0MHFR7:RWH_8P#RHRONRFHlLMHN0FDMNR0HMCsoCRP8HHs8CR0IHEFSL0JERkHF0CRM0NRM8sNClHCM8skRF00bk#
3R-a-RERH#ObFlFMMC0HR8PCH8#ER0CHR8PCH8MR8,NL,R$ER0CHR8PFH#sL,R,FR0RFbs8CkORC0ERFJk0MHC0MRN8CRslMNH83Cs
R--mHb0FDMNDR$,0RECsNClHCM8skRF00bkRlOFbCk0#ER0CFRl8kkD#-3
--
-RCaERo#HMVRFRC0ERlsCN8HMCHsR#ER0CHR#oFMRVER0CRRqHkMb0-3
-ERaCHR#oFMRVER0CFRl8kkD##RHRC0ERo#HMVRFRC0ERHARM0bk3-
--------------------------------------------------------------------------------------------------S


LDHs$NsR Q  k;
#QCR 3  #_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFHkO_Mo#HM3C8N;DD
Ck#RCHCC03#8F_Do_HON0sHED3ND
;
CHM007$RWH_8P#RH
CSoMHCsOS5
SIN_HE80SuR:ma1QQSe :c=4;S
SLH_I8S0ERm:u1QQae: S=
g;SOS0_8lFC:SRhzqa)RqpSj:=;S
Ss_CllCF8Rq:haqz)p=S:4S
S2S;
b0Fs5S
SNSRSSH:RM0R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;SRSLS:SSRRHM#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;S
SJ0kFH0CMSF:Rk#0R0D8_FOoH_OPC05FsNH_I8-0E4FR8IFM0R;j2
sSSCHlNMs8CSF:Rk#0R0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R;j2
8SSH8PHC$_L_:jSR0FkR8#0_oDFHSO
S
2;CRM878W_H;PR
s
NO0EHCkO0ssCR0FDRVWR7_P8HRRH#
-
-R0QMCNsMDHR#oDMNRO8CDNNs0MHF#H
#oDMNRsbNN,l4RFJk0J,RkHF0C_M0.R#,0bClR#:R0D8_FOoH_OPC0RFs5_RNI0H8ERR-4FR8IFM0R2jR;H
#oDMNRsbNN,l.R8lFDRR:#_08DHFoOC_POs0FRL5R_8IH0-ERR84RF0IMFRRj2
;R
R--wOkM0MHFRR0FoRC00RECJ0kFH0CMR8NMRlsCN8HMCRs31VEH0k/#Ls#0NRO0MRFMs0C#FMsHoDRNoHFs0RElHH#RlCbDl0CMCS8

MVkOF0HMHR8PRR5NRR:#_08DHFoOC_POs0F5_RNI0H8ERR-4FR8IFM0R2jR;RRL:0R#8F_Do_HOP0COFRs5LH_I8R0E-RR48MFI0jFRR22RR0sCkRsM#_08DHFoOC_POs0F;V

k0MOHRFM8RHP5RRN:0R#8F_Do_HOP0COFRs5NH_I8R0E-RR48MFI0jFRRR2;LRR:#_08DHFoOC_POs0F5_RLI0H8ERR-4FR8IFM0R2jRRs2RCs0kM0R#8F_Do_HOP0COFHsR#P

NNsHLRDC#Rkl:0R#8F_Do_HOP0COFRs5LH_I8R0E8MFI0jFRR
2;PHNsNCLDRP8HHM8C8RR:#_08DHFoOC_POs0FRN5R_8IH0-ERR84RF0IMFRRj2P;
NNsHLRDCs_ClNk8[#:0RR8#0_oDFHPO_CFO0sRR5LH_I8R0E8MFI0jFRR
2;PHNsNCLDRl0CbR_L:0R#8F_Do_HOP0COFRs5LH_I8R0E8MFI0jFRR
2;PHNsNCLDRbNb_:LRR8#0_oDFHPO_CFO0sRR5LH_I8R0E8MFI0jFRR
2;PHNsNCLDRlsC8RR:#_08DHFoOC_POs0F5IL_HE80R4-RRI8FMR0Fj;R2RL

CMoH
k
#l=R:RF5R0sEC#>R=R''jR
2;8HHP88CMRR:=N#;
kjl52=R:RNN5_8IH0-ERR;42
P8HHM8C8=R:RP8HHM8C8N5R_8IH0-ERR8.RF0IMFRRj2RR&';j'
bNb_:LR=jR''RR&R;LR
l0CbR_L:M=RFN05bLb_2+RRR''4;k
#l=R:Rl#kR0+RC_lbL8;
H8PHC5M8j:2R=FRM0RR5#5klLH_I820ER
2;VRFsHMRHR0jRFRR5NH_I8R0E-RR.2FRDFSb
H5VRRl#k5IL_HE802RR='R4'2ER0CSM
Sl0CbR_L:'=Rj&'RR
L;S#CDCS
S0bCl_:LR=FRM0b5Nb2_LRRR+';4'
MSC8VRH;#
Sk:lR=kR#l_5LI0H8ERR-4FR8IFM0R2jRR'&Rj
';Sl#k5Rj2:8=RH8PHC5M8RIN_HE80R4-RR
2;SP8HHM8C8=R:RP8HHM8C8N5R_8IH0-ERR8.RF0IMFRRj2RR&';j'
kS#l=R:Rl#kR0+RC_lbLS;
8HHP88CM5Rj2:M=RF50RRl#k5IL_HE802;R2
8CMRFDFbH;
VRR5#5klLH_I820ER'=R42'RRC0EMs
SCNl_8#[k0=R:Rl#kR5+RR''jRL&RR
2;CCD#
CSsl8_N[0k#RR:=#;kl
8CMR;HV
lsC8=R:RlsC_[N8k5#0RIL_HE80R4-RRI8FMR0Fj;R2
0sCkRsM5HR8PCH8M&8RRlsC8;R2SC

M88RH
P;
oLCH
M
-m-Rkk0b0#RN#MHol0CM
s
bF#OC#RR5L
R2LHCoMH
SVRR5LRR=j02RE
CMSHS8PCH8__L$j=R<R''4;C
SD
#CSHS8PCH8__L$j=R<R''j;C
SMH8RVC;
Mb8RsCFO#R#;R
R
-Q-RMs0CMRND#MHoNNDR#o#HMMlC0b

sCFO#5#RR2NR
oLCHSM
H5VRR_0OlCF8R4=RR02RE
CMSVSHRN5R5IN_HE80R4-R2RR='R4'2ER0CSM
SNSbs4NlRR<=M5F0N+2RR''4;S
SCCD#
SSSbNNsl<4R=;RN
CSSMH8RVS;
CCD#
bSSNlsN4=R<R
N;S8CMR;HV
8CMRFbsO#C#;b

sCFO#5#RLL2
CMoH
VSHR05ROF_l8=CRR24RRC0EMS
SH5VRRLL5_8IH0-ERR24RR'=R42'RRC0EMS
SSsbNNRl.<M=RFL052RR+4S;
S#CDCS
SSsbNNRl.<L=R;S
SCRM8H
V;S#CDCS
SbNNsl<.R=;RL
MSC8VRH;M
C8sRbF#OC#
;

FbsO#C#Rb5RNlsN4b,RNlsN.
R2PHNsNCLDRFJk0F_l8:DRR8#0_oDFHPO_CFO0sRR55IN_HE80RL+R_8IH0RE2-RR48MFI0jFRRR2;
oLCH
MSSFJk0F_l8:DR=HR8Pb5RNlsN4b,RNlsN.;R2
kSJF<0R=kRJFl0_F58DR_5NI0H8ERR+LH_I820ERR-48MFI0LFR_8IH02ER;l
SFR8D<J=Rk_F0lDF85_RLI0H8ERR-4FR8IFM0R2jR;M
C8sRbF#OC#
;
J0kFH0CM_R.#<M=RFJ05k2F0R'+R4
';
s
bF#OC#RR5J0kF,kRJFC0HM.0_#N,R,RRL2C
Lo
HMSRHV5NR55IN_HE80R4-RRG2RFLsR5IL_HE80R4-RRR22=4R''RR20MEC
0SSCRlb<J=RkHF0C_M0.R#;
DSC#SC
Sl0Cb=R<RFJk0
;RS8CMR;HV
8CMRFbsO#C#;


-m-Rkk0b0#RN#MHol0CM
s
bF#OC#RR5NRR,Ll,RFR8D2PS
NNsHLRDC0bCl4RR:#_08DHFoOC_POs0FRL5R_8IH0-ERR84RF0IMFRRj2R:=50RFE#CsRR=>'R4'2P;
NNsHLRDC0bCl.RR:#_08DHFoOC_POs0FRN5R_8IH0-ERR84RF0IMFRRj2P;
NNsHLRDC0bCl.R_j:0R#8F_Do_HOP0COF5sRRIN_HE80R.-RRI8FMR0Fj:R2=RR5FC0Es=#R>jR'';R2
sPNHDNLCCR0lRbd:0R#8F_Do_HOP0COF5sRR84RF0IMFRRj2L;
CMoHR0
SCdlbRR:=N_5NI0H8ERR-4&2RRLL5_8IH0-ERR;42R0
SC.lbRR:='R4'&CR0l_b.jS;
H5VRRlsC_8lFCRR=4RR20MEC
HSSVRR5LRR=jRR20MEC
SSSsNClHCM8s=R<RRN5LH_I8R0E-RR48MFI0jFRR
2;SDSC#RHV5OR0_8lFCRR=4MRN8RRL=CR0lRb4NRM8NRR=0bCl.RR20MECSS
SSlsCN8HMC<sR=CR0l;b4
CSSDV#HR05ROF_l8=CRRN4RM58RR8lFD=R/R2jRR8NMRNN5_8IH0-ERR24RR'=R42'RRC0EMS
SSlsCN8HMC<sR=FRM0F5l8RD2+4R''S;
S#CDCS
SSlsCN8HMC<sR=FRl8
D;SMSC8VRH;
SRS#CDH5VRR_0OlCF8R4=RR02RE
CMSHSSVRR5LRR=jRR20MEC
SSSSlsCN8HMC<sR=5RNRIL_HE80R4-RRI8FMR0Fj;R2
SSSCHD#VRR5LRR=0bCl4MRN8RRN=CR0lRb.2ER0CSM
SsSSCHlNMs8CRR<=0bCl4S;
SDSC#SC
SOSSNR#C5CR0lRbd2#RHRS
SSISSERCM""jjR
=>SSSSSlsCN8HMC<sR=FRl8SD;RS
SS
SSSSSSSCIEMjR"4="R>S
SSHSSVRR5lDF8RR/=jRR20MEC
SSSSsSSCHlNMs8CRR<=LRR+lDF8;S
SSCSSD
#CSSSSSCSslMNH8RCs<l=RF;8D
SSSSMSC8VRH;S
SSSS
SSSSIMECRj"4">R=
SSSSVSHRl5RFR8D/j=RR02RESCMRSR
SSSSSlsCN8HMC<sR=RRL-FRl8
D;SSSSS#CDCS
SSSSSsNClHCM8s=R<R8lFDS;
SSSSCRM8H
V;SSSSSS
SSISSERCM""44R
=>SSSSSRHV5FRl8/DR=RRj2ER0CSM
SSSSSlsCN8HMC<sR=FRM0F5l8RD2+4R''S;
SSSSCCD#
SSSSsSSCHlNMs8CRR<=lDF8;S
SSCSSMH8RVS;
SSSS
SSSSESICFMR0sEC#>R=
SSSSkSMD
D;SSSSCRM8OCN#;S
SS8CMR;HV
CSSD
#CSHSSVRR5LRR=jRR20MEC
SSSSlsCN8HMC<sR=5RNRIL_HE80R4-RRI8FMR0Fj;R2
SSSCCD#
SSSSlsCN8HMC<sR=FRl8
D;SCSSMH8RVS;
S8CMR;HV
CS
Mb8RsCFO#
#;
R--mbk0kN0R#o#HMMlC0b

sCFO#5#RR,NRRRL,0bCl,kRJF20RRN
PsLHND0CRC4lbR#:R0D8_FOoH_OPC0RFs5_RLI0H8ERR-4FR8IFM0R2jR:5=RREF0CRs#='>R42'R;N
PsLHND0CRC.lbR#:R0D8_FOoH_OPC0RFs5_RNI0H8ERR-4FR8IFM0R2jR;N
PsLHND0CRC.lb_:jRR8#0_oDFHPO_CFO0sRR5NH_I8R0E-RR.8MFI0jFRR:2R=RR5FC0Es=#R>jR'';R2
sPNHDNLCCR0lRbd:0R#8F_Do_HOP0COF5sRRIN_HE80R4-RRI8FMR0Fj;R2
sPNHDNLCCR0l_bd4RR:#_08DHFoOC_POs0FRN5R_8IH0-ERR8.RF0IMFRRj2=R:RF5R0sEC#>R=R''4R
2;PHNsNCLDRl0Cb:cRR8#0_oDFHPO_CFO0sRR5NH_I8R0E-RR48MFI0jFRR=2:RF5R0sEC#>R=R''4R
2;
oLCH
MRSl0Cb:.R=4R''RR&0bCl.;_j
CS0lRbd:'=Rj&'RRl0Cb4d_;H
SVRR5L=R/R2jRRC0EMS
SOCN#R05ROF_l82CRR
H#SISSERCM4>R=
SSSH5VRR=LRRl0CbN4RMN8RR0=RC.lbR02RE
CMSSSSJ0kFH0CMRR<=0bCldS;
SDSC#SC
SJSSkHF0CRM0<0=RC;lb
SSSCRM8H
V;S
SSSISSERCMj>R=
SSSJ0kFH0CMRR<=J0kF;S
SSS
SSCIEM0RFE#CsR
=>SMSSk;DD
SSS
CSSMO8RN;#C
DSC#SC
S#ONCRR50lO_FR8C2#RH
SSSIMECR=4R>S
SSRHV55RNNH_I8R0E-RR42RR='R4'2ER0CSM
SJSSkHF0CRM0<0=RC.lb;S
SS#CDCS
SSkSJFC0HM<0R=CR0l;bdRS
SS8CMR;HVSSR
SSS
SESICjMRR
=>SJSSkHF0CRM0<0=RCclb;SR
SSS
SESICFMR0sEC#>R=
SSSMDkD;S
SCRM8OCN#;C
SMH8RV
;SCRM8bOsFC;##
M
C80RsD
;
DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOs_NH30EN;DD
Ck#RCHCC03#8F_Do_HOkHM#o8MC3DND;C

M00H$QR7e#RH
RRRRMoCCOsH5R
SRIRRHE80RRR:HCM0oRCs:4=R(S;
RRRRs8IH0RER:MRH0CCos=R:R;4(
RSRRIRNHE80RH:RMo0CC:sR=;Rg
RSRRIRLHE80RH:RMo0CC:sR=2RU;R
RRFRbs
05SqRS:MRHR8#0_oDFHPO_CFO0sI5NHE80RR-48MFI0jFR2S;
SRA:H#MR0D8_FOoH_OPC05FsL8IH0-ER4FR8IFM0R;j2
7SSQ7eQ RR:FRk0#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
)SS Qvqh:7SR0FkR8#0_oDFHPO_CFO0sI5sHE80-84RF0IMF2Rj2C;
M78RQ
e;
s
NO0EHCkO0sOCRC_DDDCCPDVRFRe7QR
H#
FSOlMbFCRM078W_HSP
oCCMs5HO
NSS_8IH0RES:1umQeaQ S;
SIL_HE80SuR:ma1QQ;e 
0SSOF_l8RCS:ahqzp)qRS;
SlsC_8lFChR:q)azqSp
S
2;SsbF0S5
SSNRSRS:H#MR0D8_FOoH_OPC05FsNH_I8-0E4FR8IFM0R;j2
LSSRSSS:MRHR8#0_oDFHPO_CFO0s_5LI0H8ER-48MFI0jFR2S;
SFJk0MHC0RS:FRk0#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;S
SsNClHCM8sRS:FRk0#_08DHFoOC_POs0F5IL_HE80-84RF0IMF2Rj;S
S8HHP8LC_$S_j:kRF00R#8F_Do
HOS;S2
MSC8FROlMbFC;M0
C
Lo
HM
VSH_MoCC0sNCD_bkR#:H5VRN8IH0>ER=IRLHE802CRoMNCs0SC
So#HMRNDNk_NG:RRR8#0_oDFHPO_CFO0sI5NHE80RI8FMR0FjR2;RS
S#MHoNLDR_GNkRRR:#_08DHFoOC_POs0F5HLI8R0E8MFI0jFR2R;R
#SSHNoMD_RJNRkGR#:R0D8_FOoH_OPC05FsN8IH08ERF0IMF2Rj;
RRSHS#oDMNRNs_kRGR:0R#8F_Do_HOP0COFLs5I0H8EFR8IFM0R;j2RSR
LHCoMS
SNk_NG=R<R""jRq&R;S
SLk_NG=R<R""jRA&R;

SSkSlD:04RWR7_P8H
SSSoCCMsRHOlRNb5S
SS_SNI0H8E>R=RHNI8+0E4S,
SLSS_8IH0=ER>IRLHE80+
4,SSSS0lO_FR8C=j>R,S
SSCSslF_l8=CR>
R4S2SS
SSSb0FsRblNRS5
SNSSRR=>qk_NGS,
SLSSRR=>Lk_NGS,
SJSSkHF0CRM0=J>R_GNk,S
SSCSslMNH8RCs=s>R_GNk
SSS2
;

SRSS_HVoCCMsCN0_R4:H5VRs8IH0>ERRHLI820ERMoCC0sNCS
SS S)vhqQ7=R<RhBmea_17m_pt_QBea Bmj)5,IRsHE80RL-RI0H8ERR2&_RsN5kGL8IH0-ER4FR8IFM0R;j2
SSSCRM8oCCMsCN0R_HVoCCMsCN0_
4;
SRSS_HVoCCMsCN0_R.:H5VRs8IH0<ER=IRLHE802CRoMNCs0SC
S)SS Qvqh<7R=_RsN5kGs8IH04E-RI8FMR0Fj
2;SCSSMo8RCsMCNR0CHoV_CsMCN_0C.
;
RSSSHoV_CsMCN_0CdH:RVIR5HE80RN>RI0H8Eo2RCsMCN
0CSSSS7QQe7< R=mRBh1e_ap7_mBtQ_Be a5m)jI,RHE80RN-RI0H8ERR2&_RJN5kGN8IH0-ERR84RF0IMF2Rj;S
SS8CMRMoCC0sNCVRH_MoCC0sNC;_d
S
RSVSH_MoCC0sNC:_cRRHV58IH0<ER=IRNHE802CRoMNCs0SC
S7SSQ7eQ =R<RNJ_kIG5HE80-84RF0IMF2Rj;S
SS8CMRMoCC0sNCVRH_MoCC0sNC;_c
MSC8CRoMNCs0HCRVC_oMNCs0bC_D;k#
SS
HoV_CsMCN_0ClkHM#H:RVNR5I0H8ERR<L8IH0RE2oCCMsCN0
#SSHNoMD_RNNRkGR#:R0D8_FOoH_OPC05FsL8IH08ERF0IMF2Rj;
RRSHS#oDMNRNL_kRGR:0R#8F_Do_HOP0COFLs5I0H8EFR8IFM0R;j2RSR
So#HMRNDJk_NG:RRR8#0_oDFHPO_CFO0sI5LHE80RI8FMR0FjR2;RS
S#MHoNsDR_GNkRRR:#_08DHFoOC_POs0F5HLI8R0E8MFI0jFR2R;R
CSLo
HMS_SNNRkG<B=Rm_he1_a7pQmtB _eB)am5Rj,L8IH0-ERRHNI8R0E+2R4Rq&R;S
SLk_NG=R<RhBmea_17m_pt_QBea Bmj)5,2R4RA&R;

SSkSlD:04RWR7_P8H
SSSoCCMsRHOlRNb5S
SS_SNI0H8E>R=RHLI8+0E4S,
SLSS_8IH0=ER>IRLHE80+
4,SSSS0lO_FR8C=j>R,S
SSCSslF_l8=CR>
R4S2SS
SSSb0FsRblNRS5
SNSSRR=>Nk_NGS,
SLSSRR=>Lk_NGS,
SJSSkHF0CRM0=J>R_GNk,S
SSCSslMNH8RCs=s>R_GNk
SSS2
;

SRSS_HVoCCMsCN0_R4:H5VRs8IH0>ERRHLI820ERMoCC0sNCS
SS S)vhqQ7=R<RhBmea_17m_pt_QBea Bmj)5,IRsHE80RL-RI0H8ERR2&_RsN5kGL8IH0-ERR84RF0IMF2Rj;S
SS8CMRMoCC0sNCVRH_MoCC0sNC;_4
S
RSVSH_MoCC0sNC:_.RRHV5HsI8R0E<L=RI0H8Eo2RCsMCN
0CSSSS)q vQRh7<s=R_GNk5HsI8-0E4FR8IFM0R;j2
SSSCRM8oCCMsCN0R_HVoCCMsCN0_
.;
SRSS_HVoCCMsCN0_Rd:H5VRI0H8ERR>L8IH0RE2oCCMsCN0
SSSSe7QQR7 <B=Rm_he1_a7pQmtB _eB)am5Rj,I0H8ERR-L8IH02ERRJ&R_GNk5HLI8R0E-RR48MFI0jFR2S;
SMSC8CRoMNCs0HCRVC_oMNCs0dC_;R

SHSSVC_oMNCs0cC_:VRHRH5I8R0E<L=RI0H8Eo2RCsMCN
0CSSSS7QQe7< R=_RJN5kGI0H8ER-48MFI0jFR2S;
SMSC8CRoMNCs0HCRVC_oMNCs0cC_;C
SMo8RCsMCNR0CHoV_CsMCN_0ClkHM#
;
CRM8ODCD_PDCC
D;
