@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Wa_QBh_]tqh 
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
V`H8RCVm_ep1)]q B7_m
7 
sRRCIoRHFM8IRR=j
;
RDRNI#N$RR@@5#bFCC8oR	OD2CRLo
HMRRRRH5VR`pme_1)  1a_Qqthp=R!RL4'jL2RCMoH
RRRRHRRV!R5I8HMF&IR&0R#N_s0CMPC0=R=RL4'4R2
RRRRRIRRHFM8I=R<RL4'4R;
RRRRR#CDCVRHRH5IMI8FRR&&C_M8CMPC0=R=RL4'4R2
RRRRRIRRHFM8I=R<RL4'jR;
RCRRMR8
RCRRDR#CLHCoMR
RRRRRI8HMF<IR='R4L
j;RRRRC
M8RMRC8`

CHM8V/R/Rpme_q1])_ 7B m7
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 aQ_Wh]_Bq ht_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R#R500Ns_CCPM&0R&IR!HFM8Iy2Ryf4R#L0ND0C5C_#0CsGb24r*:Rf9|R->!8CM_CCPM
0;RMRC8Fbsb0Cs$`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRsRbFsbC0q$R1)1 aQ_Wh]_Bq ht__XZm1h_aaq)_  ehua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R!H5IMI8F2-R|>!R55#fHkMM	F5IM#s0N0P_CC2M02
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_hWQ_qB]h_t XmZ_h _a1 a_X_u)uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RH5IMI8F2-R|>!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Wa_QBh_]tqh Z_X__mh _h7 he a;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRI8HMFRI2|R->5f!5HM#k	IMFMM5C8P_CC2M02
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)aW_QhBh]qtu _:#RN#0CsRFbsb0Cs$qR51)1 aQ_Wh]_Bq ht_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFR#ENR0MFRNOEM8oCRDPNkLCRCsVFCHRIMI8FRRH#O#DFC28";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 aQ_Wh]_Bq ht__XZm1h_aaq)_  ehua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aW_QhBh]qtX _Zh_m_q1a) a_ea h_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#s0N0P_CCRM0O0FMN#HMRFXRs"RZ2R;
RRRRRqRR_1q1 _)aW_QhBh]qtX _Zh_m_1a aX_ uu)_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aW_QhBh]qtX _Zh_m_1a aX_ uu)_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RRRRRqRR_1q1 _)aW_QhBh]qtX _Zh_m_7 h_  ehua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aW_QhBh]qtX _Zh_m_7 h_  ehua_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5M"C8P_CCRM0O0FMN#HMRFXRs"RZ2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRv1_q1a )_hWQ_qB]h_t uN:R#l#kCsRbFsbC05$Rq 11)Wa_QBh_]tqh 2_u;


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqv_1)1 aQ_Wh]_Bq ht__XZm1h_aaq)_  ehua_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aW_QhBh]qtX _Zh_m_q1a) a_ea h_;u2
RRRRRRRRqv_1)1 aQ_Wh]_Bq ht__XZmah_ _1a )Xu_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_Wh]_Bq ht__XZmah_ _1a )Xu_;u2
RRRRRRRRqv_1)1 aQ_Wh]_Bq ht__XZm h_h 7_ea h_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_Wh]_Bq ht__XZm h_h 7_ea h_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_ho

CsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_CsI8HMFFI_b:CM
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRRRRRN#0sC0_P0CMRR&&!MIH82FIRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8_FIFMbCRPOFC8sC"
2;
RRRRORRFsPC_MIH8:FI
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52R`pme_1)  1a_Qqthp=R!RL4'j02REksFokEF0R
RRRRRRRRRRRRRRRRRR5RR5N#0sC0_P0CMRR&&!MIH82FIR4yy
RRRRRRRRRRRRRRRRRRRR!R5C_M8CMPC0&R&RMIH82FIRjr*:Rf9y
y4RRRRRRRRRRRRRRRRRRRRRM5C8P_CCRM0&I&RHFM8IR222R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05I8HMFOIRFsPCC28";R
RRCRRM/8R/#LNHOORFsPCN
oCRRRRC
M8
8CMoCCMsCN0
M`C8RHV/m/ReBp_m)e _
mh
