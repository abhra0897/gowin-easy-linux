@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)aa_Q"v ;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"

V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
RMRHHN0HDCRLo
HMRRRRH5VR~N55OF0HMM_F_IMC_N#0s=0R=mR`eQp_t)hm  _hWa_1q2)aR
||RRRRRRRRRNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqa|2R|R
RRRRRRRRR50NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)a2L2RCMoH
RRRRFRRPCD_sssF_"05QCDDoRNDPkNDCCR#0FRVsNRbsCNl0RCsNHO0FFM_MC_MI0_#N"s02R;
RCRRMR8
R8CM
H
`VV8CRpme_q1])_ 7B m7RR

RosCRMIH8RFI=;Rj
HRRMo0CCHsRRj=R;R

RINDNR$#@5@RbCF#8RoCO2D	RoLCHRM
RHRRV`R5m_ep)  1aQ_1tphqRR!=4j'L2CRLo
HMRRRRRVRHRI5!HFM8I&R&RN#0sC0_P0CMRR==44'L2CRLo
HMRRRRRRRRI8HMF<IR='R4L
4;RRRRRRRRH=R<RlMk_#O	;R
RRRRRC
M8RRRRRDRC#HCRVIR5HFM8IL2RCMoH
RRRRRRRRRHV5=HR=RR4&5&RNHO0FFM_MC_MI0_#NRs0!`=Rm_ep)  1ah_m_Wh _q1a)|aR|R
RRRRRRRRRRRRRRRRRRRRRRN#0sC0_P0CMRR!=44'L2R2
RRRRRRRRRMIH8RFI<4=R';Lj
R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)R
&&RRRRRRRRRRRR#s0N0P_CCRM0=4=R'2L4
RRRRRRRRHRRRR<=M_klO;	#
RRRRRRRR#CDCVRHRR5H!4=R2R
RRRRRRRRRH=R<R-HRR
4;RRRRRMRC8/R/RRHV5MIH82FI
RRRR8CM
RRRR#CDCCRLo
HMRRRRRHRIMI8FRR<=4j'L;R
RRRRRH=R<R
j;RRRRC
M8RMRC8`

CHM8V/R/Rpme_q1])_ 7B m7
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 aQ_avu _;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5N#0sC0_P0CMRR&&!MIH82FIR>|=RC50#C0_G2bsrk*Ml	_O#
9;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_vaQ  _)1_ am1h_aaq)_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R#R500Ns_CCPMR02|R=>5RR
RRRRRRRRRRRRRRRRRRRRR055C_#0CsGb2Mr*kOl_	2#9
RSRRRRRRRRRRRRRF
sRRRRRRRRRRRRRRRRRRRRRR5R500C#_bCGs*2rjk:Ml	_O#9-4R4yyRN#0sC0_P0CM2SR
RRRRRRRRRRRR2R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aa Qv_) )__mh1)aqa;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
IRRHFM8I-R|>#R!00Ns_CCPM
0;RMRC8Fbsb0Cs$


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
bRRsCFbsR0$q 11)aa_Q_v XmZ_ha_1q_)auR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RI!5HFM8I|2R-5>R!H5f#	kMMMFI5N#0sC0_P0CM2;22
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 aQ_avX _Zh_m_Wh _q1a)ua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5MIH82FIR>|-R55!fkH#MF	MI#M500Ns_CCPM2022R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aa Qv__XZmah_ _1a )Xu_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RIR5HFM8I|2R-5>R!H5f#	kMMMFI5#0C0G_Cb2s22R;
R8CMbbsFC$s0
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
oRRCsMCN
0CRRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_ep)  1ah_m_Wh _q1a)
a2RRRRRRRRR_Rqq 11)aa_Q_v uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_vaQ 2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRRH#MRF0a )zR0IHERHM#ObCHCVH8kRMl	_O#$ROO#DCRFVslER0C0R#N_s0CMPC0;"2
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_1)  ma_h _hWa_1q2)a
RRRRRRRRqRR_1q1 _)aa Qv_1)  ma_ha_1q_)auR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_vaQ  _)1_ am1h_aaq)_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHM#RFa0R)Rz IEH0H#MRbHCOV8HCRlMk_#O	ROO$DRC#VlsFRC0ERN#0sC0_P0CM"
2;RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0=`=Rm_ep m)))h_m_Wh _q1a)
a2RRRRRRRRR_Rqq 11)aa_Q_v  _))m1h_aaq)_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 aQ_av  _)m)_ha_1q_)auR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0Q5"DoDCN#DR00NsRCCPMI0REEHOR#ENRFsCOsOkCL8RCsVFCFROlCbD0MHFRRFVOsksCRM0I8HMF2I";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 aQ_avX _Zh_m_q1a)ua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aa Qv__XZm1h_aaq)_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#s0N0P_CCRM0O0FMN#HMRFXRs"RZ2R;
RRRRRHRRVNR5OF0HMM_F_IMC_N#0s!0R=mR`eQp_t)hm  _hWa_1q2)a
RRRRRRRRqRR_1q1 _)aa Qv__XZmhh_ 1W_aaq)_
u:RRRRRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aa Qv__XZmhh_ 1W_aaq)_
u2RRRRRRRRRRRRCCD#RDFP_sCsF0s_50"#N_s0CMPC0FROMH0NMX#RRRFsZ;"2
RRRRRRRRqq_1)1 aQ_avX _Zh_m_1a aX_ uu)_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aa Qv__XZmah_ _1a )Xu_
u2RRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
R
RRRRRC
M8RRRRRmR`eqp_1v1z RR:LHCoMRR:F_PDNk##lRC
RRRRRHRRVNR5OF0HMM_F_IMC_N#0s!0R=mR`e)p_ a1 __mhh_ W1)aqaR2
RRRRRRRRRqv_1)1 aQ_avu _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aa Qv_;u2
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_1)  ma_h _hWa_1q2)a
RRRRRRRRvRR_1q1 _)aa Qv_1)  ma_ha_1q_)auR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_vaQ  _)1_ am1h_aaq)_;u2
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)a
RRRRRRRRvRR_1q1 _)aa Qv_) )__mh1)aqa:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)aa_Q_v  _))m1h_aaq)_;u2
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )_vaQ Z_X__mh1)aqa:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)aa_Q_v XmZ_ha_1q_)au
2;RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_epQmth)h _ 1W_aaq)2R
RRRRRRRRRv1_q1a )_vaQ Z_X__mhh_ W1)aqa:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_vaQ Z_X__mhh_ W1)aqa2_u;R
RRRRRR_Rvq 11)aa_Q_v XmZ_h _a1 a_X_u)uR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_vaQ Z_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R

RRRRR8CM
RRRR`RRm_epQmth): RRoLCH:MRRDFP_MHoF
sCRRRRRRRR/8/RFFRM0MEHo
R;RRRRRMRC8R
RRRRR8NCVkRD0RRRR:MRHHN0HDPRFDs_Cs_Fs0"5"2R;
RCRRMN8O#RC
R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
H
RVOR5FsPCN_oCDCCPD=R!Re`mpm_Be_ )h mh2CRLoRHM:PRFDF_OP
CsRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RFROP_CsI8HMFFI_b:CM
RRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRR#RR00Ns_CCPM&0R&IR!HFM8I22R
RRRRRRRRRRRRRRRRFRRPOD_FsPC_"05I8HMFFI_bRCMOCFPs"C82
;
RORRFsPC_MIH8_FIO#DFCR:
RFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRMIH8RFI&5&RH=R=R&4R&NR5OF0HMM_F_IMC_N#0s!0R=mR`e)p_ a1 __mhh_ W1)aqa|R|RN#0sC0_P0CMRR!=44'L2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2
RRRRRRRRRRRRRRRRR
R2RRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05I8HMFOI_DCF#RPOFC8sC"
2;RMRC8/R/LHN#OFROPNCso
C
RVRHRe5mpm_Be_ )Bhm) m)_hL2RCMoHRF:RPOD_FsPC_sOFM
CsRHRRVNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqaL2RCMoHRF:RPOD_FsPC_MIH8_FIsCC#0R#
R
RRRRRROCFPsH_IMI8F_#sCC:0#
RRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRRRRRRRRRRRRRRN#0sC0_P0CMRR&&I8HMFRI22R
RRRRRRRRRRRRRRRRRRDFP_POFC0s_5H"IMI8F_#sCCR0#OCFPs"C82R;
RMRC8R
RCRM8/F/OssMCRPOFCosNCR

CRM8/e/mpm_Be_ )h mh
M
C8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



