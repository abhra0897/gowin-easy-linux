-- $Header: //synplicity/mapacx/mappers/xilinx/lib/gen_virtex5/cmp_eq.vhd#1 $
@EH
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;C

M00H$JRC_CCDl0CMR
H#RRRRb0Fs5,NjR,LjR,N4R,L4R,N.R,L.RHD0MRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRR00Fk:kRF00R#8F_Do2HO;M
C8JRC_CCDl0CM;


NEsOHO0C0CksRMCJRRFVCCJ_DCClMH0R##
SHNoMD4R0R#:R0D8_FOoH;

SSlOFbCFMMv0RzYXB_Rp
SFSbs50R
RRRSpSSmRR:FRk0#_08DHFoOR;
RSRSSRBQ:MRHR8#0_oDFH
O;RSRRSQS7RH:RM0R#8F_Do;HO
RRRS1SSRH:RM0R#8F_Do
HOR2SS;C
SMO8RFFlbM0CM;-
S-0N0skHL0LCRD	NO_GLFRRFVvBzXYRR:ObFlFMMC0#RHRk0sCL;
CMoH
4S0RR<=5RN.GsMFR2L.R8NMR45NRFGMs4RL2MRN8NR5jMRGFLsRj
2;RRRRl_kGH0M#Rv:RzYXB_Rp
RRRRRbRRFRs0l5Nb1>R=R,04RR
RRRRRRmRpRR=>Dk0F0R,
RRRRRBRRQ>R=RHD0MR,
RRRRR7RRQ>R=R''j2C;
MC8RJ
M;
H
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;C

M00H$JRC_CCDl0CM_F0IL#H0R
H#RRRRb0Fs5,NjR,LjR,N4R,L4RHD0MRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRR00Fk:kRF00R#8F_Do2HO;M
C8JRC_CCDl0CM_F0IL#H0;


NEsOHO0C0CksRMCJRRFVCCJ_DCClM00_IHFL0H#R##
SHNoMD4R0R#:R0D8_FOoH;

SSlOFbCFMMv0RzYXB_Rp
SFSbs50R
RRRSpSSmRR:FRk0#_08DHFoOR;
RSRSSRBQ:MRHR8#0_oDFH
O;RSRRSQS7RH:RM0R#8F_Do;HO
RRRS1SSRH:RM0R#8F_Do
HOR2SS;C
SMO8RFFlbM0CM;-
S-0N0skHL0LCRD	NO_GLFRRFVvBzXYRR:ObFlFMMC0#RHRk0sCL;
CMoH
4S0RR<=5RN4GsMFR2L4R8NMRj5NRFGMsjRL2R;
RlRRkHG_MR#0:zRvX_BYpR
RRRRRRFRbsl0RN1b5RR=>0R4,
RRRRRRRRRpm=D>R00Fk,R
RRRRRRQRBRR=>DM0H,R
RRRRRRQR7RR=>'2j';M
C8JRCM
;

LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
M
C0$H0R_CJClDCC_M0FLMCHH0R#R
RRFRbsN05jL,RjD,R0RHM:MRHR8#0_oDFH
O;RRRRRRRRRRRRRFD0kR0:FRk0#_08DHFoO
2;CRM8CCJ_DCClMF0_MHCL0
;

ONsECH0Os0kCJRCMVRFR_CJClDCC_M0FLMCHH0R##
SHNoMD4R0R#:R0D8_FOoH;

SSlOFbCFMMv0RzYXB_Rp
SFSbs50R
RRRSpSSmRR:FRk0#_08DHFoOR;
RSRSSRBQ:MRHR8#0_oDFH
O;RSRRSQS7RH:RM0R#8F_Do;HO
RRRS1SSRH:RM0R#8F_Do
HOR2SS;C
SMO8RFFlbM0CM;-
S-0N0skHL0LCRD	NO_GLFRRFVvBzXYRR:ObFlFMMC0#RHRk0sCL;
CMoH
4S0RR<=5RNjGsMFR2Lj;R
RRkRlGM_H#:0RRXvzBpY_
RRRRRRRRsbF0NRlbR51=0>R4
,RRRRRRRRRp=mR>0RDF,k0
RRRRRRRRRBQ=D>R0,HM
RRRRRRRRR7Q='>Rj;'2
8CMRMCJ;



LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
M
C0$H0RuBv_R THR#
RoRRCsMCHIO5HE80RH:RMo0CC:sR=;42
RRRRsbF0:5qRRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRR:RARRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRRTR RF:Rk#0R0D8_FOoH2C;
MB8Rv u_T
;

ONsECH0Os0kCCRODDD_CDPCRRFVB_vu HTR#V

k0MOHRFMVOkM_sCsFCs5JH_I8R0E:MRH0CCoss2RCs0kM0R#soHMR
H#LHCoMR
RH5VR5_CJI0H8E=R>R262RC0EMR
RRCRs0Mks52"";R
RCCD#
RRRR0sCk5sM"sCsF2s";R
RCRM8H
V;CRM8VOkM_sCsF
s;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FOVRC_DDDCCPDRR:NEsOHO0C0CksRRH#VOkM_sCsFIs5HE802
;
SMOF#M0N00RHC0sNHRFM:MRH0CCos=R:RH5I820E/
d;SMOF#M0N0CRslMNH8RCs:MRH0CCos=R:RH5I820ER8lFR
d;RRRR#MHoN8DRN_0N0Rlb:0R#8F_Do_HOP0COF5sRI0H8ERR-4FR8IFM0R;j2
R
RRFROlMbFCRM0CCJ_DCClMH0R#R
RRRRRRFRbsN05jL,RjN,R4L,R4N,R.L,R.D,R0:HMRRHM#_08DHFoOR;
RRRRRRRRRRRRRRRRDk0F0RR:FRk0#_08DHFoO
2;RRRRCRM8ObFlFMMC0
;
RRRRObFlFMMC0JRC_CCDl0CM_F0IL#H0R
H#RRRRRRRRb0Fs5,NjR,LjR,N4R,L4RHD0MH:RM0R#8F_Do;HO
RRRRRRRRRRRRRRRR0RDFRk0:kRF00R#8F_Do2HO;R
RRMRC8FROlMbFC;M0
O
SFFlbM0CMR_CJClDCC_M0FLMCHH0R#R
RRRRRRFRbsN05jL,RjD,R0:HMRRHM#_08DHFoOR;
RRRRRRRRRRRRRRRRDk0F0RR:FRk0#_08DHFoO
2;RRRRCRM8ObFlFMMC0L;
CMoH
jSzRH:RVI5RHE80R4>R2CRoMNCs0SC
LHCoMR
RRjRz4RR:CCJ_DCClMR0
RRRRRRRRRRRRRbRRFRs0l5Nb
RSSRRNj=q>R5,j2RR
RRRRRRRRRRRRRRRRRL=jR>5RAj
2,SRSRN=4R>5Rq4R2,
RRRRRRRRRRRRRRRRLRR4>R=R4A52S,
SNRR.>R=R.q52
,RRRRRRRRRRRRRRRRRR.RLRR=>A25.,R
RRRRRRRRRRRRRR0RDH=MR>4R''R,
RRRRRRRRRRRRRDRR00FkRR=>8NN0_b0l52j2;C
SMo8RCsMCN;0C
R
RRRRRRSR
z:4RR5HVR8IH0=ERRR42oCCMsCN0
CSLo
HMSTS RR<=q25jRFGMs5RAj
2;S8CMRMoCC0sNC
;
RRRRz:.RRsVFR0LH_8HMCHGRMRR405FRHs0CNF0HMRR-4R2RoCCMsCN0
RRRRRRRRoLCHRM
RRRRRRRRRzRR.:4RR_CJClDCC
M0RRRRRRRRRRRRRRRRb0FsRblN5S
SN=jR>5RqdH*L0M_H82CG,RR
RRRRRRRRRRRRRLRRj>R=RdA5*0LH_8HMC,G2
NSS4>R=Rdq5*0LH_8HMC+GRR,42RR
RRRRRRRRRRRRRR4RLRR=>A*5dL_H0HCM8GRR+4
2,S.SNRR=>q*5dL_H0HCM8GRR+.R2,
RRRRRRRRRRRRRRRRRL.=A>R5Ld*HH0_MG8CR.+R2R,
RRRRRRRRRRRRRDRR0RHM=8>RN_0N05lbL_H0HCM8GRR-4
2,RRRRRRRRRRRRRRRRDk0F0>R=R08NNl_0bH5L0M_H82CG2R;
RRRRRCRRMo8RCsMCN;0C
z
Sd:qRR5HVRlsCN8HMC=sRRN.RMI8RHE80R4>R2CRoMNCs0SC
LHCoMS
SzRd4:JRC_CCDl0CM_F0IL#H0
SSSb0FsRblN5S
SSjSNRR=>qH5I8R0E-,.2
SSSSRLj=A>R58IH0-ERR,.2
SSSSRN4=q>R58IH0-ER4
2,SSSSL=4R>5RAI0H8ERR-4
2,SSSSDM0HR8=>N_0N05lbHs0CNF0HMRR-4
2,SSSSDk0F0>R=R2 T;C
SMo8RCsMCN;0C
z
SdRR:HRV5sNClHCM8sRR=4MRN8HRI8R0E>2R4RMoCC0sNCL
SCMoH
zSSd:4RR_CJClDCC_M0FLMCHS0
SFSbsl0RN
b5SSSSN=jR>5RqI0H8E4R-2S,
SLSSj>R=RIA5HE80R4-R2S,
SDSS0RHM=N>800N_lHb50NCs0MHFR4-R2S,
SDSS00FkRR=> ;T2
MSC8CRoMNCs0
C;
RRRRRRRRz
ScRR:HsV5CHlNMs8CRj=RR8NMR8IH0RER>2R4RMoCC0sNCL
SCMoH
RRRRTS RR<=8NN0_b0l5CH0sHN0F-MRR;42RS

CRM8oCCMsCN0;C

MR8RODCD_PDCC
D;
