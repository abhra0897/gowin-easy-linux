@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)wa_Q_wmQ h7X
";
HR`MkOD8"CR#_08F_PD0	N#3
E"R`R
HCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0M`C
CHM8V/R/m_epQahQ_tv1
R
RH0MHHRNDLHCoMR
RRVRHRC58b=0E=
j2RRRRRDFP_sCsF0s_5D"QDNCoDNRPDRkCVRFsbNNslCC0sCR8bR0EIOEHEkRl#L0RCCR#0FR0RDPNkoCRs0CNC0sRERNMj;"2
CRRM
8
`8HVCmVRe1p_] q)7m_B7
 
R0HMCsoCR0OM;H
RMHH0NODRM=0RR
j;
NRRD$IN#@R@5#bFCC8oR	OD2CRLo
HMRRRRRVRHRm5`e)p_ a1 _t1QhRqp!4=R'2LjRoLCHRM
RRRRRHRRV{R5bEk#!,=jb!Fb=Rj}=.=R'jL42CRLoRHM/b/Rk
#ERRRRRRRRRVRHRO55M+0RR#bkE<2R=CR8b20ERoLCHRM
RRRRRRRRRORRM<0R=MRO0RR+bEk#;R
RRRRRRRRRC
M8RRRRRRRRC
M8RRRRRRRRCCD#RRHV5k{b#=E!jF,bbj!=}=R=RL.'jR42LHCoM/R/RbbF
RRRRRRRRHRRVOR5M>0R=FRbbL2RCMoH
RRRRRRRRRRRR0OMRR<=ORM0-FRbbR;
RRRRRRRRR8CM
RRRRRRRR8CM
RRRRRRRR#CDCVRHRb5{k!#E=bj,F=b!j=}R='R.L244RoLCH/MR/kRb#&ERRbbF
RRRRRRRRHRRV!R5#kHlDM0NC#Fk_#bkEF_bbL2RCMoH
RRRRRRRRRRRRQ//ptp qupRzR1]qRh7u
muRRRRRRRRRMRC8R
RRRRRRRRRCCD#RoLCHRM
RRRRRRRRRHRRV5R5ORM0+kRb#-ERRbbF2RR>80CbEL2RCMoH
RRRRRRRRRRRR/RR/ me)mwpWR"
RRRRRRRRRCRRMR8
RRRRRRRRRCRRDR#CH5VR50OMRb+Rk2#ERb<RFRb2LHCoMR
RRRRRRRRRRRRR/h/z7w )p
mWRRRRRRRRRRRRC
M8RRRRRRRRRRRRCCD#RoLCHRM
RRRRRRRRRRRRR0OMRR<=ORM0+kRb#-ERRbbF;R
RRRRRRRRRRMRC8R
RRRRRRRRRC
M8RRRRRRRRC
M8RRRRRMRC8R
RRRRRCCD#RoLCHRM
RRRRRORRM<0R=;Rj
RRRRCRRMR8
R8CM
C
`MV8HRR//m_ep1)]q B7_m
7 
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_wwQmh_Q7_ Xm)e wWpm_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RkRb#&ER&5R!!l#HkND0MkCF#k_b#bE_F&bR&kRb#&ER&FRbb|2R-5>R50OMRb+RkR#E-FRbb<2R=CR8b20E;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)wa_Q_wmQ h7Xh_z7w )p_mWuR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RF5bb&R&R!!5#kHlDM0NC#Fk_#bkEF_bb&R&R#bkE&R&RbbF2&R&Rk5b#=ER=RRj|5|R5M5O0RR+bEk#Rb-RFRb2<8=RCEb02222R>|-RO55M+0RR#bkE>2R=FRbb
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_wwQmh_Q7_ XQ ppt_qpu]z1_uum_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R!bEk#RR&&b2Fb;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_wwQmh_Q7_ XXmZ_hz_u1u]_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5HM#k	IMFMk5b#2E22R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)awmQw_7Qh XX_Zh_m_uum_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R!R55#fHkMM	F5IMb2Fb2
2;RMRC8Fbsb0Cs$R

RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##s
0
RRRRRRRRq1_q1a )_wwQmh_Q7_ Xm)e wWpm_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)awmQw_7Qh mX_ew )p_mWuR2
RRRRRCRRDR#CF_PDCFsss5_0"VwHFPRFCDsVF8IRCO0C0"C82
;
RRRRRRRRq1_q1a )_wwQmh_Q7_ Xz h7)mwpW:_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_wwQmh_Q7_ Xz h7)mwpW2_u
RRRRRRRR#CDCPRFDs_Cs_Fs0w5"HRVFkCM8sFVDICR800COC28";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 aQ_wwQm_hX7 __XZmuh_z_1]uR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_Q_wmQ h7XZ_X__mhu]z1_
u2RRRRRRRRCCD#RDFP_sCsF0s_5k"b#OERFNM0HRM#XsRFR2Z";R

RRRRRqRR_1q1 _)awmQw_7Qh XX_Zh_m_uum_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)awmQw_7Qh XX_Zh_m_uum_
u2RRRRRRRRCCD#RDFP_sCsF0s_5F"bbFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
R
RRRRRRVRHR#5!HDlk0CNMF_k#bEk#_bbF2CRLoRHM:_RNNC##sV0_H_VFHCM8GD_HDNCoDk_b#bE_FRb
RRRRRRRRRqq_1)1 aQ_wwQm_hX7 _pQp ptq_1uz]m_uu:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_Q_wmQ h7Xp_Qpq tpz_u1u]_muu_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5D"QDNCoDHR#l0kDNFMCkb#RkR#EbRFb8CC0O80C"
2;RRRRRRRRC
M8RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
R
RRRRRR_Rvq 11)wa_Q_wmQ h7Xe_m p)wmuW_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_wwQm_hX7 _ me)mwpW2_u;R

RRRRRvRR_1q1 _)awmQw_7Qh zX_h)7 wWpm_
u:RRRRRRRRNk##lbCRsCFbsR0$51q1 _)awmQw_7Qh zX_h)7 wWpm_;u2
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )_wwQmh_Q7_ XXmZ_hz_u1u]_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_wwQm_hX7 __XZmuh_z_1]u
2;
RRRRRRRRqv_1)1 aQ_wwQm_hX7 __XZmuh_muu_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_wwQm_hX7 __XZmuh_muu_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRH5VR!l#HkND0MkCF#k_b#bE_FRb2LHCoMRR:l#_N#0Cs_VVHFM_H8_CGHCDDo_NDbEk#_bbF
RRRRRRRRvRR_1q1 _)awmQw_7Qh QX_ptp qup_z_1]u_muuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_wwQmh_Q7_ XQ ppt_qpu]z1_uum_;u2
RRRRRRRR8CM
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_ho

CsMCN
0C
VRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRHV5pme_eBm A)_qB1Q_2mhRoLCH:MRRDFP_POFCLs_NO#H
RRR
RRROCFPsH_VVbF_k:#E
RRROCFPssRbFsbC05$RR5@@bCF#8RoCO2D	R`55m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRbRRkR#E&b&RF=bR=2Rj2R
RRRRRF_PDOCFPs5_0"VVHFk_b#OERFsPCC28";R

RFROP_CsVFHV_bbF:R
RRPOFCbsRsCFbsR0$5@R@5#bFCC8oR	OD25R5`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRbRFb&b&RkR#E=j=R2R2
RRRRRDFP_POFC0s_5H"VVbF_FObRFsPCC28";R
RCRM8/N/L#RHOOCFPsCNo
R
RH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR

RFROP_CsVFHV_DVkDR:
RFROPRCsbbsFC$s0R@5R@F5b#oC8CDRO	52R5e`mp _)1_ a1hQtq!pR='R4LRj2&
&RRRRRR/R/R#ONCERICRsCF$MDR#bkE#RHRk0sCMRN8HRVVoFRFRC#0VFRk
DDRRRRR5R55#bkE=R!j&2R&OR5M+0RbEk#RR==80CbE&2R&bR5F=bR=2j2RR||
R
RRRRR/O/RNR#CIEH0Rl#HkND0MkCF#kRb#NERMb8RFNbRMV8RHRVFo#FCRR0FVDkD
RRRR5RR5bbFRR!=j&2R&bR5kR#E!j=R2&R&RO55M-0RRbbFRb+Rk2#ERR==80CbE&2R&RR
RRRRRH5#l0kDNFMCkb#_k_#Eb2Fb2R2
RRRRR22R
RRRRDFP_POFC0s_5H"VVVF_kRDDOCFPs"C82
;
RORRFsPC_VVHFl_Cb:0$
RRROCFPssRbFsbC05$RR5@@bCF#8RoCO2D	R`55m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRR/RR/NRO#ICRECCsRDFM$FRbb#RHRk0sCMRN8HRVVoFRFRC#0CFRl$b0
RRRR5RR5F5bb=R!RRj2&5&RbEk#RR==j&2R&5R5ORM0-FRbb=2R=2Rj2|R|RR

RRRRRR//OCN#R0IHEHR#l0kDNFMCkb#RkR#ENRM8bRFbNRM8VFHVRCoF#FR0RbCl0R$
RRRRRb55F!bR=2RjRR&&5#bkE=R!RRj2&5&R50OMRb-RF+bRR#bkE=2R=2RjRR&&
RRRR5RR#kHlDM0NC#Fk_#bkEF_bb222
RRRR2RRRR2
RRRRRDFP_POFC0s_5H"VVCF_l$b0RPOFC8sC"
2;
RRROCFPsH_VV#F_HDlk0CNMF_k#bEk#_bbF:R
RRPOFCbsRsCFbsR0$5@R@5#bFCC8oR	OD25R5`pme_1)  1a_Qqthp=R!RL4'j&2R&kRb#&ER&FRbb
22RRRRRPRFDF_OP_Cs0V5"H_VF#kHlDM0NC#Fk_#bkEF_bbFROPCCs8;"2
CRRM/8R/sOFMRCsOCFPsCNo
C
RM/8R/pme_eBm h)_m
h 
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m
