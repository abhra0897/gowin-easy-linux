
@ER--=========m==F=FF=========================================FmFF========-
-RR=RB$FbsEHo0BR52jR.4.c-jR46tHFIMCR1lFHOMO8k0RFsaECOMFFDoB$RFp3,0
83-=-RRRRRRRRRRRRRRRRRRRRRRDqDRosHER0#sCC#s8PC3-
-R====================================================================-=
--
-R_R_RRRRR_R_RRRRR_R_
R--R\\RRRRR/\RRRRRR/RR/RwRrHRDCMCNlR9RRRHbsl$_#ME3P8-
-R\RRRR\R/\R/RR\R/RR/RrRR7OC#s0HbHRFM9]Re7VpRk0MOHNFMD$R#MC0E#RH#DsHLN
s$-R-RRRR\\//RRRR\\//RRRRRRHral0C#NRlbRRR9WRC8qRko.4nR6j:j:Rdj.6j4
R--RRRR\/RRRRRR\/RRRRRRRPRrCHs#FRMRR9RRR.433-4
-RRRR\RR/RRRR\RR/RRRRRRR

---=-R=========F=mF=F=========================================mFFF========
-

-------------------------N-bOo	NCDRoFDLN-----------------------------
-
p)QAqR)YHCCC;zR
1H RC3CC#_08DHFoO4_4nNc3DRD;
Ck#R Q  a317m_pt_QBqa)Q]p3qpk;
#QCR 3  1_a7pQmtBh_z1hQt q73p
p;
Buqi qtRlOFbCFMMR0#Q
1RRNRR0H0sLCk0RM#$_NLDOL	_FRG:LDFFCRNM;R
RR0N0skHL0#CR$LM_D	NO_GLFRRFVBbFlFMMC0:#RRObN	CNoRRH#0Csk;R
RR0N0skHL0LCRD	NO_GLF_8bN_MbH:0R#soHM;R
RR0N0skHL0#CR$MM_FkbsM:CRRFLFDMCN;R
RR0N0skHL0GCRON_lb#:R0MsHoR;
R0RN0LsHkR0CGlO_NFbRVFRBlMbFC#M0Rb:RNNO	oHCR#DR"k;0"R-S
-ObN	CNoRLoDR
H#-#-SHNoMD1Rt):hRR8#0_oDFH:OR=4R''-;
-8CMRLoD;-
-b	NONRoCL$F8RLoDR-
-CRM8o;DL
----------------------------t--1-)--------------------------------------B

mmvuha hR)t1RR
RRmRu)5aR
RRRRRRRR1Rt):QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR)t1RB:RFFlbM0CMRRH#0Csk;-
-------------------------p4za-----------------------------B-
mmvuha hRapz4RR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXj2"R;R
RRmRu)5aR
wSRRF:Rk#0R0D8_FOoH;R
RRRRRRQRRjRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh a
;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRa4:FRBlMbFCRM0H0#Rs;kC
0N0skHL0GCRON_lbVRFRapz4RR:ObFlFMMC0#RHRk"D0
";S-
-------------------------p.zaR----------------------------B-
mmvuha hRapz.RR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXj2"R;R
RRmRu)5aR
RRRSRRw:kRF00R#8F_Do;HO
RRRSjRQRH:RM0R#8F_Do;HO
RRRS4RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRa.:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:.RRlOFbCFMMH0R#DR"k;0"
------------------------p--z-ad-----------------------------m
Bvhum RhapdzaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"j2"R;R
RRmRu)5aR
RRRSRRw:kRF00R#8F_Do;HO
RRRSjRQRH:RM0R#8F_Do;HO
RRRS4RQRH:RM0R#8F_Do;HO
RRRS.RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:dRRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapzdRR:ObFlFMMC0#RHRk"D0
";-------------------------z-pa-cR----------------------------
vBmu mhhpaRzRac
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"jjRj"2R;
RuRRmR)a5R
RRwSRRF:Rk#0R0D8_FOoH;R
RRQSRjRR:H#MR0D8_FOoH;R
RRQSR4RR:H#MR0D8_FOoH;R
RRQSR.RR:H#MR0D8_FOoH;R
RRQSRdRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRac:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:cRRlOFbCFMMH0R#DR"k;0"
------------------------p--zRa6-----------------------------m
Bvhum Rhap6zaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"jjjjj"jjR
2;RRRRuam)RR5
RRRSwRR:FRk0#_08DHFoOR;
RRRSQ:jRRRHM#_08DHFoOR;
RRRSQ:4RRRHM#_08DHFoOR;
RRRSQ:.RRRHM#_08DHFoOR;
RRRSQ:dRRRHM#_08DHFoOR;
RRRSQ:cRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVp6zaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRa6:FROlMbFCRM0H"#RD"k0;-
-------------------------pnzaR----------------------------
-
Bumvmhh azRpa
nRRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjj2"R;R
RRmRu)5aR
RRRSRRw:kRF00R#8F_Do;HO
RRRSjRQRH:RM0R#8F_Do;HO
RRRS4RQRH:RM0R#8F_Do;HO
RRRS.RQRH:RM0R#8F_Do;HO
RRRSdRQRH:RM0R#8F_Do;HO
RRRScRQRH:RM0R#8F_Do;HO
RRRS6RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:nRRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapznRR:ObFlFMMC0#RHRk"D0
";-------------------------z-pa-(R----------------------------
m
Bvhum Rhap(zaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR
2;RRRRuam)RR5
RRRSwRR:FRk0#_08DHFoOR;
RRRSQ:jRRRHM#_08DHFoOR;
RRRSQ:4RRRHM#_08DHFoOR;
RRRSQ:.RRRHM#_08DHFoOR;
RRRSQ:dRRRHM#_08DHFoOR;
RRRSQ:cRRRHM#_08DHFoOR;
RSRRRRQ6:MRHR8#0_oDFH
O;RSRRRRQn:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRapz(RR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVp(zaRO:RFFlbM0CMRRH#"0Dk"-;
-------------------------apzU-R--------------------------
--
vBmu mhhpaRzRaU
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"2R;
RuRRmR)a5R
RRwSRRF:Rk#0R0D8_FOoH;R
RRQSRjRR:H#MR0D8_FOoH;R
RRQSR4RR:H#MR0D8_FOoH;R
RRQSR.RR:H#MR0D8_FOoH;R
RRQSRdRR:H#MR0D8_FOoH;R
RRQSRcRR:H#MR0D8_FOoH;R
RRQSR6RR:H#MR0D8_FOoH;R
RRQSRnRR:H#MR0D8_FOoH;R
RRQSR(RR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRaU:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:URRlOFbCFMMH0R#DR"k;0"
------------------------v--z-X.-----------------------------B

mmvuha hRXvz.RR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;SjR1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzRX.:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.p6za-----------------------------
-
Bumvmhh azRvXp._zRa6
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_pa:6RRlBFbCFMMH0R#sR0k
C;-------------------------z-vXp._z-an-----------------------------B

mmvuha hRXvz.z_pa
nRRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apznRR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvz.z_pa-(-----------------------------
m
Bvhum Rhav.zX_apz(RR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;SjR1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.p(zaRB:RFFlbM0CMRRH#0Csk;-
-------------------------v.zX_apzU----------------------------
--
vBmu mhhvaRz_X.pUzaRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRaU:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.vUzX-----------------------------
-
Bumvmhh azRvXv._zRXU
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_vX:URRlBFbCFMMH0R#sR0k
C;-------------------------z-vXv._znX4-----------------------------
-
Bumvmhh azRvXv._znX4RR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXv._znX4RB:RFFlbM0CMRRH#0Csk;-
-------------------------v.zX_Xvzd-.-----------------------------
m
Bvhum Rhav.zX_Xvzd
.RRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_Xvzd:.RRlBFbCFMMH0R#sR0k
C;-------------------------z-vX-c-----------------------------
m
Bvhum RhavczXRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RRQ.:MRHR8#0_oDFHRO;
QSRdRR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
RR14:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvX:cRRlBFbCFMMH0R#sR0k
C;-------------------------z-vX-U-----------------------------
m
Bvhum RhavUzXRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RRQ.:MRHR8#0_oDFHRO;
QSRdRR:H#MR0D8_FOoH;R
SQ:cRRRHM#_08DHFoOS;
RRQ6:MRHR8#0_oDFH
O;SnRQRH:RM0R#8F_Do;HO
QSR(RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
RR14:MRHR8#0_oDFH
O;S.R1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzRXU:FRBlMbFCRM0H0#Rs;kC
------------------------v--znX4-----------------------------B

mmvuha hRXvz4RnR
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
SQ:.RRRHM#_08DHFoO
;RSdRQRH:RM0R#8F_Do;HO
QSRcRR:H#MR0D8_FOoH;R
SQ:6RRRHM#_08DHFoOS;
RRQn:MRHR8#0_oDFH
O;S(RQRH:RM0R#8F_Do;HO
QSRURR:H#MR0D8_FOoH;R
SQ:gRRRHM#_08DHFoOS;
RjQ4RH:RM0R#8F_Do;HO
QSR4:4RRRHM#_08DHFoOS;
R.Q4RH:RM0R#8F_Do;HO
QSR4:dRRRHM#_08DHFoOS;
RcQ4RH:RM0R#8F_Do;HO
QSR4:6RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;S4R1RH:RM0R#8F_Do;HO
1SR.RR:H#MR0D8_FOoH;R
S1:dRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz4:nRRlBFbCFMMH0R#sR0k
C;-------------------------z-vX-d.----------------------------
m
Bvhum RhavdzX.
RRRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
QSR.RR:H#MR0D8_FOoH;SR
RRQd:MRHR8#0_oDFH
O;ScRQRH:RM0R#8F_Do;HO
QSR6RR:H#MR0D8_FOoH;R
SQ:nRRRHM#_08DHFoOS;
RRQ(:MRHR8#0_oDFH
O;SURQRH:RM0R#8F_Do;HO
QSRgRR:H#MR0D8_FOoH;R
SQR4j:MRHR8#0_oDFH
O;S4RQ4RR:H#MR0D8_FOoH;R
SQR4.:MRHR8#0_oDFH
O;S4RQdRR:H#MR0D8_FOoH;R
SQR4c:MRHR8#0_oDFH
O;S4RQ6RR:H#MR0D8_FOoH;R
SQR4n:MRHR8#0_oDFH
O;S4RQ(RR:H#MR0D8_FOoH;R
SQR4U:MRHR8#0_oDFH
O;S4RQgRR:H#MR0D8_FOoH;R
SQR.j:MRHR8#0_oDFH
O;S.RQ4RR:H#MR0D8_FOoH;R
SQR..:MRHR8#0_oDFH
O;S.RQdR:RH#MR0D8_FOoH;R
SQR.c:MRHR8#0_oDFH
O;S.RQ6RR:H#MR0D8_FOoH;R
SQR.n:MRHR8#0_oDFH
O;S.RQ(RR:H#MR0D8_FOoH;R
SQR.U:MRHR8#0_oDFH
O;S.RQgRR:H#MR0D8_FOoH;R
SQRdj:MRHR8#0_oDFH
O;SdRQ4RR:H#MR0D8_FOoH;SR
RR1j:MRHR8#0_oDFH
O;S4R1RH:RM0R#8F_Do;HO
1SR.RR:H#MR0D8_FOoH;R
S1:dRRRHM#_08DHFoOS;
RR1c:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXRd.:FRBlMbFCRM0H0#Rs;kC
------------------------q--p-z------------------------------B

mmvuha hRzqpRR
RR RthQ )BRR5RR
RRRRRRqRR7:7RRaQh )t RR:=j
R;RRRRRSRRRA1zRQ:Rhta  :)R=RR4;R
RRRRRRqRR7z71ARR:Q hatR ):.=RRR;
RRRRRRRSh: RRaQh )t RR:=d
R;RRRRRSRRRRt :hRQa  t)=R:R;cR
pSR RR:Q hatR ):6=R;R
RRRRRRBSRz:uRRaQh )t RR:=n
R;RRRRRRRRRhB7RQ:Rhta  :)R=RR(;R
RRRRRRBRRz7uBhRR:Q hatR ):U=R;R
SvazpRQ:Rhta  :)R=;Rg
qSRpvz_mR7 :hRQa  t)=R:RRj
R2RR;RS
RuRRmR)a5R
S1Rzv:zRma0R#8F_Do;HO
BSRmRza:zRma0R#8F_Do;HOSR
SQ:jRRRQh#_08DHFoOS;
R:Q4RRQh#_08DHFoOS;
R:QdRRQh#_08DHFoOS;
RhBQ:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRqzRR:BbFlFMMC0#RHRk0sC-;
-------------------------7--w-wR-----------------------------B

mmvuha hRw7wRR
RR RthQ )BRR5QahQRL:RH:0R=jR''S2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw:wRRlBFbCFMMH0R#sR0k
C;-------------------------7--wRw ---------------------------------B

mmvuha hRw7w RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S RBRQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w: RRlBFbCFMMH0R#sR0k
C;-------------------------w7w1-R------------------------------
--
vBmu mhh7aRwRw1
RRRRht  B)QRQ5Rh:QaR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
1SR :aRRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV71wwRB:RFFlbM0CMRRH#0Csk;-
--------------------------w-7w-1 -------------------------------------B

mmvuha hRw7w1
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
1SR :aRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV71ww RR:BbFlFMMC0#RHRk0sC-;
---------------------7--wRw)---------------------------------
-
Bumvmhh awR7w
)RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
)SR a1 RQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:)RRlBFbCFMMH0R#sR0k
C;-------------------------7--w w)R------------------------------------
-
Bumvmhh awR7wR) 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S)  1aRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw w)RB:RFFlbM0CMRRH#0Csk;-
--------------------------w-7w-u--------------------------------------B

mmvuha hRw7wuRR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S)Ru a1 :hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wuRR:BbFlFMMC0#RHRk0sC-;
-------------------------w7wu- R--------------------------------------------
m
Bvhum Rha7uww RR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S)Ru a1 RQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRu :FRBlMbFCRM0H0#Rs;kC
----------------------------w-7w-BR-----------------------------
--
vBmu mhh7aRwRwB
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRwB:FRBlMbFCRM0H0#Rs;kC
----------------------------w-7wRB -----------------------------------------
--
vBmu mhh7aRw wBRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R Bpq:)RRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Bww RR:BbFlFMMC0#RHRk0sC-;
-------------------------w7wh-R-----------------------------
m
Bvhum Rha7hwwRR
RR RthQ )BRR5QahQRL:RH:0R=jR''S2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRwh:FRBlMbFCRM0H0#Rs;kC
----------------7--w whR--------------------------------
-
Bumvmhh awR7wRh 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SB: RRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww RR:BbFlFMMC0#RHRk0sC-;
------------------------7hww1-R------------------------------
--
vBmu mhh7aRw1whRR
RR RthQ )BRR5QahQ:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S1R a:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:1RRlBFbCFMMH0R#sR0k
C;----------------------------7hww1- -------------------------------------
m
Bvhum Rha7hww1
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
1SR :aRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww1: RRlBFbCFMMH0R#sR0k
C;-----------------------------w7wh-)---------------------------------
m
Bvhum Rha7hww)RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R)1R a:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:)RRlBFbCFMMH0R#sR0k
C;-------------------------7--w)wh -R----------------------------------
--
vBmu mhh7aRw)wh RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R)1R a:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whR) :FRBlMbFCRM0H0#Rs;kC
----------------------------w7wh-u--------------------------------------B

mmvuha hRw7wh
uRRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRhu:FRBlMbFCRM0H0#Rs;kC
------------------------7--wuwh -R------------------------------------------
--
vBmu mhh7aRwuwh RR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S)Ru a1 RQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w huRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--wBwhR--------------------------------------------B

mmvuha hRw7wh
BRRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRhB:FRBlMbFCRM0H0#Rs;kC
----------------------------w-7w hBR-------------------------------------------
m
Bvhum Rha7hwwB
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w hBRB:RFFlbM0CMRRH#0Csk;-
------------------------------p-7R----------------------------------------
--
vBmu mhh7aRpRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRR:BbFlFMMC0#RHRk0sC-;
------------------------7-p ---------------------------------
-
Bumvmhh apR7 RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp: RRlBFbCFMMH0R#sR0k
C;-----------------------------B7pR------------------------------------B

mmvuha hRB7pRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R Bpq:)RRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7BRR:BbFlFMMC0#RHRk0sC-;
----------------------------7 pBR------------------------------------B

mmvuha hRB7p RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRB :FRBlMbFCRM0H0#Rs;kC
----------------------------p-7u-R----------------------------------
-
Bumvmhh apR7uRR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;SS
RRt:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rpu:FRBlMbFCRM0H0#Rs;kC
----------------------------p-7u- R---------------------------------
--
vBmu mhh7aRpRu 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
Su1)  :aRRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7u: RRlBFbCFMMH0R#sR0k
C;------------------------7Rph-----------------------------------------
-
Bumvmhh apR7hRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:hRRlBFbCFMMH0R#sR0k
C;-----------------------------h7p -----------------------------------
m
Bvhum Rha7 phRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7h: RRlBFbCFMMH0R#sR0k
C;-----------------------------h7pB-R----------------------------------
-
Bumvmhh apR7h
BRRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7BphRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--p hBR------------------------------------B

mmvuha hRh7pB
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Bph RR:BbFlFMMC0#RHRk0sC-;
----------------------------7uphR------------------------------------B

mmvuha hRh7puRR
RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;SS
RRt:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7uphRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--p huR------------------------------------B

mmvuha hRh7pu
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7pu: RRlBFbCFMMH0R#sR0k
C;---------------------A-Qz-w----------------------------------
--
vBmu mhhQaRARzw
RRRR)uma
R5RRRRSRRm:zRma0R#8F_Do;HO
RRRRQSRRQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVARQz:wRRlBFbCFMMH0R#sR0k
C;-----------------------------A-mz-w--------------------------------------B

mmvuha hRzmAwRR
RuRRmR)a5R
RRRRSmRR:mRza#_08DHFoOR;
RSRRR:QRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVmwAzRB:RFFlbM0CMRRH#0Csk;-
----------------------------------A-az-w--------------------------B

mmvuha hRzaAwRR
RuRRmR)a5R
RRRRSmRR:mRza#_08DHFoOR;
RSRRR:QRRRQh#_08DHFoOR;
RSRRRRm :hRQR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzaAwRR:BbFlFMMC0#RHRk0sC-;
-------------------------Q--mwAz--------------------------------
m
Bvhum RhaQzmAwRR
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSQ:mRRmQhz#aR0D8_FOoH;R
RRSRRRRQR:hRQRRRR#_08DHFoOS;
RRm :hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQzmAwRR:BbFlFMMC0#RHRk0sC-;
--------------------------------Q)77)------------------------
--
vBmu mhhQaR7)7)RR
RR RthQ )B
R5S_TjQahQRL:RH:0R=jR''S;
TQ4_hRQa:HRL0=R:R''j
RRRRS2;
RRRR)uma
R5SjRTRm:Rz#aR0D8_FOoH;R
ST:4RRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
)SR a1 :hRQR8#0_oDFHSO;
BSRpRi:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ)77)RR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRV7RQ7R)):FRBlMbFCRM0H"#RTRj,T;4"
--------------------------------7-Q7-)1-------------------------
-
Bumvmhh a7RQ7R)1
RRRRht  B)QRS5
TQj_hRQa:HRL0=R:R''4;T
S4h_QQ:aRR0LHRR:='
4'RRRR2
;SRRRRuam)RS5
RRTj:zRma0R#8F_Do;HO
TSR4RR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S R1aQ:Rh0R#8F_Do;HOSR
SB:piRRQh#_08DHFoOS;
R:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7Q7):1RRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFQVR717)RB:RFFlbM0CMRRH#",TjR"T4;-
------------------------------Q--7B7)-------------------------
--
vBmu mhhQaR7B7)RR
RR RthQ )BRR5
jST_QQhaRR:LRH0:'=Rj
';S_T4QahQRL:RH:0R=jR''R
RR;R2SR
RRmRu)5aR
TSRjRR:mRza#_08DHFoOS;
RRT4:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )Q:Rh0R#8F_Do;HOSR
SB:piRRQh#_08DHFoOS;
R:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7Q7):BRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFQVR7B7)RB:RFFlbM0CMRRH#",TjR"T4;-
------------------------------Q--7u7)-------------------------
--
vBmu mhhQaR7u7)RR
RR RthQ )BRR5
jST_QQhaRR:LRH0:'=R4
';S_T4QahQRL:RH:0R=4R''R
RR;R2SR
RRmRu)5aR
TSRjRR:mRza#_08DHFoOS;
RRT4:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
Su1)  Ra:Q#hR0D8_FOoH;SS
RiBp:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ7R)u:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVQ)77uRR:BbFlFMMC0#RHRj"T,4RT"-;
-------------------------Q--7_7)v- v---------------------------------
--
vBmu mhhQaR7_7)vR v
 SthQ )B
R5S1St)R h:FRLFNDCM=R:RDVN#
C;S1Sp)R hRL:RFCFDN:MR=sR0kSC
2S;
uam)RS5
SRTj:kRF00R#8F_Do;HOSS
ST:4RR0FkR8#0_oDFHSO;
7SSRH:RM0R#8F_Do;HO
BSS RR:H#MR0D8_FOoH;S
SQiBpRH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SqSW7j7)RH:RM0R#8F_Do;HO
RSRRqSW747)RH:RM0R#8F_Do;HO
RSRRqSW7.7)RH:RM0R#8F_Do;HO
)SSq)77jRR:H#MR0D8_FOoH;R
SR)RSq)774RR:H#MR0D8_FOoH;R
SR)RSq)77.RR:H#MR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ)77_vv RB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7Q7) _vvRR:BbFlFMMC0#RHRj"T,4RT"-;
-----------------------------7-m7-))---------------------B

mmvuha hR7m7)
)RRRRRt  h)RQB5mRBhq1ahQaRhRQa:0R#8F_DoRHO:'=Rj2'R;RS
RuRRmR)a5SR
R:TRRamzR8#0_oDFHSO;
7SRjRR:Q#hR0D8_FOoH;R
S7:4RRRQh#_08DHFoOS;
RRB :hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOS;
R1)  :aRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7m7):)RRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFmVR7)7)RB:RFFlbM0CMRRH#",7jR"74;-
------------------------------7m7)-1---------------------
m
Bvhum Rham)771RR
RtRR )h Q5BRRhBm1haqahRQQ:aRR8#0_oDFH:OR=4R'';R2SR
RRmRu)5aRRR
STRR:mRza#_08DHFoO
;SSjR7RQ:Rh0R#8F_Do;HO
7SR4RR:Q#hR0D8_FOoH;R
SB: RRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH;R
S1R a:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7R)1:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVm)771RR:BbFlFMMC0#RHRj"7,4R7"-;
-----------------------------7-m7-)B---------------------B

mmvuha hR7m7)
BRRRRRt  h)RQB5mRBhq1ahQaRhRQa:0R#8F_DoRHO:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSjR7RQ:Rh0R#8F_Do;HO
7SR4Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFH
O;S RBRH:RM0R#8F_Do;HO
BSRp) q:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7R)B:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVm)77BRR:BbFlFMMC0#RHRj"7,4R7"-;
-----------------------------7-m7-)u---------------------B

mmvuha hR7m7)
uRRRRRt  h)RQB5mRBhq1ahQaRhRQa:0R#8F_DoRHO:'=R42'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSjR7RQ:Rh0R#8F_Do;HO
7SR4Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFH
O;S RBRH:RM0R#8F_Do;HO
uSR)  1aQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR7u7)RB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7m7):uRRlBFbCFMMH0R#7R"j7,R4
";----------------------------m)77_vv ------------------------------------
m
Bvhum Rham)77_vv RR
RR RthQ )BS5
S)t1 :hRRFLFDMCNRR:=V#NDCS;
S)p1 RhR:FRLFNDCM=R:Rk0sCR
RR;R2
RRRR)uma
R5STSRjRR:FRk0#_08DHFoO
;SSTSR4RR:FRk0#_08DHFoO
;SSaSRBRpi:MRHR8#0_oDFH
O;SuSRBRpi:MRHR8#0_oDFH
O;SBSR RR:H#MR0D8_FOoH;S
SR1)  :aRRRHM#_08DHFoOS;
SjR7RH:RM0R#8F_Do;HO
RSS7:4RRRHM#_08DHFoOS;
SXRaRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7v)_ :vRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFmVR7_7)vR v:FRBlMbFCRM0H"#R7Rj,7;4"
----------------------------------------7-Q -1c-----------------------------
-
Bumvmhh a7RQ R1c
 SthQ )B
R5S1St): hADFFCRNM:V=RNCD#;S
Sp 1)hF:AFNDCM=R:Rk0sC2
S;u
SmR)a5S
S7RR:Q#hR0D8_FOoH;S
S)  1aRR:Q#hR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SpwBiRR:Q#hR0D8_FOoH;S
SuiBpRQ:Rh0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do;HO
TSS.RR:mRza#_08DHFoOS;
SRTd:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7c 1RB:RFFlbM0CMRRH#0Csk;-
-------------------------Q17 c _vv--------------------------------
--
vBmu mhhQaR7c 1_vv Ro
SCsMCH
O5S1St): hADFFCRNM:V=RNCD#;S
Sp 1)hF:AFNDCM=R:Rk0sC2
S;u
Sm5)a
7SS,1)  Ba, RR:Q#hR0D8_FOoH;S
SQiBp,pwBiB,up:iRRRQh#_08DHFoOS;
S7Wq7,)jW7q7)W4,q)77.RR:Q#hR0D8_FOoH;S
S)7q7))j,q)774q,)7.7)RQ:Rh0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do;HO
TSS.RR:mRza#_08DHFoOS;
SRTd:zRma0R#8F_Do
HOS;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 c _vvRR:BbFlFMMC0#RHRk0sC-;
---------------------------------Q--eCH8F-------------------------------
m
Bvhum RhaQ8eHC
FRRRRRt  h)RQB5S
SR1Rt)R h:FRLFNDCM=R:Rpwq1
 ;SRSRp 1)hRR:LDFFCRNM:a=R)
z RRRR2R;
RuRRmR)a5S
S7RR:Q#hR0D8_FOoH;R
RRBRS RR:H#MR0D8_FOoH;S
S)  1aRR:Q#hR0D8_FOoH;S
SBQqpARR:Q#hR0D8_FOoH;S
SwiBpRQ:Rh0R#8F_Do;HO
uSSBRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVReCH8FRR:BbFlFMMC0#RHRk0sC-;
---------------------------------7-Q -1U------------------------------------
m
Bvhum RhaQ17 URR
RtRR )h Q5BR
tSR1h) RA:RFCFDN:MR=NRVD;#C
pSR1h) RA:RFCFDN:MR=sR0kRC
R2RR;R
RRmRu)5aR
7SS,1)  Ba, RR:Q#hR0D8_FOoH;S
SwiBp,puBiRR:Q#hR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH;S
ST:.RRamzR8#0_oDFH
O;SdSTRm:Rz#aR0D8_FOoH;S
ST:cRRamzR8#0_oDFH
O;S6STRm:Rz#aR0D8_FOoH;S
ST:nRRamzR8#0_oDFH
O;S(STRm:Rz#aR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7U 1RB:RFFlbM0CMRRH#0Csk;-
----------------------Q--7U 1_vv ----------------------------
m
Bvhum RhaQ17 U _vvRR
RtRR )h Q5BR
tSR1h) RA:RFCFDN:MR=NRVD;#C
pSR1h) RA:RFCFDN:MR=sR0kRC
R2RR;R
RRmRu)5aR
7SS,1)  Ba, RR:Q#hR0D8_FOoH;S
SwiBp,pQBiB,up:iRRRQh#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoOS;
SRT.:zRma0R#8F_Do;HO
TSSdRR:mRza#_08DHFoOS;
SRTc:zRma0R#8F_Do;HO
TSS6RR:mRza#_08DHFoOS;
SRTn:zRma0R#8F_Do;HO
TSS(RR:mRza#_08DHFoOS;
S7Wq7R)j:MRHR8#0_oDFH
O;SqSW747)RH:RM0R#8F_Do;HO
WSSq)77.RR:H#MR0D8_FOoH;S
S)7q7):jRRRHM#_08DHFoOS;
S7)q7R)4:MRHR8#0_oDFH
O;SqS)7.7)RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ _1UvR v:FRBlMbFCRM0H0#Rs;kC
------------------------------------Q--74 1j--------------------------------
--
vBmu mhhQaR74 1jRR
RtRR )h Q5BR
tSR1h) RA:RFCFDN:MR=NRVD;#C
pSR1h) RA:RFCFDN:MR=sR0kRC
R2RR;R
RRmRu)5aR
7SS,1)  Ba, RR:Q#hR0D8_FOoH;S
SwiBp,puBiRR:Q#hR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH;S
ST:.RRamzR8#0_oDFH
O;SdSTRm:Rz#aR0D8_FOoH;S
ST:cRRamzR8#0_oDFH
O;S6STRm:Rz#aR0D8_FOoH;S
ST:nRRamzR8#0_oDFH
O;S(STRm:Rz#aR0D8_FOoH;S
ST:URRamzR8#0_oDFH
O;SgSTRm:Rz#aR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR74 1jRR:BbFlFMMC0#RHRk0sC-;
------------------------m)1 c----------------------------
--
vBmu mhhmaR1c )Rt
S )h Q5BR
tSS1h) RL:RFCFDN:MR=qRwp;1 
pSS1h) RL:RFCFDN:MR=)RazS 
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SjaXRH:RM0R#8F_Do;HO
aSSX:4RRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SBSup:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SpwBiRR:H#MR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 cRR:BbFlFMMC0#RHRk0sC-;
----------------m)1 c _vv--------------------------------B

mmvuha hR m1)vc_ 
vRSht  B)QRS5
S)t1 :hRRFLFDMCNRR:=w1qp S;
Sp]WRL:RFCFDN:MR=qRwp;1 
pSS1h) RL:RFCFDN:MR=)RazS 
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SjaXRH:RM0R#8F_Do;HO
aSSX:4RRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SBSup:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SpwBiRR:H#MR0D8_FOoH;S
SaiBpRH:RM0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR1c )_vv RB:RFFlbM0CMRRH#0Csk;-
------------------e-mHF8C---------------------------------
-
Bumvmhh aeRmHF8CRt
S )h Q
B5S1St)R h:FRLFNDCM=R:Rpwq1
 ;S1Sp)R h:FRLFNDCM=R:Rza) 2
S;u
SmR)a5S
S7:jRRRHM#_08DHFoOS;
SR74:MRHR8#0_oDFH
O;S.S7RH:RM0R#8F_Do;HO
7SSdRR:H#MR0D8_FOoH;S
S7:cRRRHM#_08DHFoOS;
SR76:MRHR8#0_oDFH
O;SnS7RH:RM0R#8F_Do;HO
BSS RR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SRST:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVReCH8FRR:BbFlFMMC0#RHRk0sC-;
-----------------m--1U )---------------------------------
--
vBmu mhhmaR1U )RR
RR RthQ )B
R5RRRRS1Rt)R h:FRLFNDCM=R:Rpwq1
 ;RRRRS1Rp)R h:FRLFNDCM=R:Rza) R
RR;R2
RRRR)uma
R5RRRRRSRR7:jRRRHM#_08DHFoOR;
RRRRR7RS4RR:H#MR0D8_FOoH;R
RRRRRR.S7RH:RM0R#8F_Do;HO
RRRRRRRSR7d:MRHR8#0_oDFH
O;RRRRRSRR7:cRRRHM#_08DHFoOR;
RRRRR6S7RH:RM0R#8F_Do;HO
RRRRRRRSR7n:MRHR8#0_oDFH
O;RRRRRSRR7:(RRRHM#_08DHFoOR;
RRRRRaRSX:jRRRHM#_08DHFoOR;
RSRRaRX4:MRHR8#0_oDFH
O;SRRRR.aXRH:RM0R#8F_Do;HO
RSRRXRadRR:H#MR0D8_FOoH;R
SRBRR RR:H#MR0D8_FOoH;RRRRR
SRuRRBRpi:MRHR8#0_oDFH
O;SRRRR1)  :aRRRHM#_08DHFoOS;
RRRRwiBpRH:RM0R#8F_Do;HO
RRRRRRRSRTj:zRma0R#8F_Do;HO
RRRRRRRSRT4:zRma0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rm R)U:FRBlMbFCRM0H0#Rs;kC
----------------1-m _)Uv- v-----------------------------
--
vBmu mhhmaR1U )_vv Rt
S )h Q
B5S1St)R h:FRLFNDCM=R:Rpwq1
 ;SWS]pRR:LDFFCRNM:w=Rq p1;S
Sp 1)hRR:LDFFCRNM:a=R)
z S
2;S)uma
R5SjS7RH:RM0R#8F_Do;HO
7SS4RR:H#MR0D8_FOoH;S
S7:.RRRHM#_08DHFoOS;
SR7d:MRHR8#0_oDFH
O;ScS7RH:RM0R#8F_Do;HO
7SS6RR:H#MR0D8_FOoH;S
S7:nRRRHM#_08DHFoOS;
SR7(:MRHR8#0_oDFH
O;SXSajRR:H#MR0D8_FOoH;S
SaRX4:MRHR8#0_oDFH
O;SXSa.RR:H#MR0D8_FOoH;S
SaRXd:MRHR8#0_oDFH
O;S SBRH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSwp:iRRRHM#_08DHFoOS;
SpaBiRR:H#MR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 U _vvRR:BbFlFMMC0#RHRk0sC-;
-----------------m--14 )j-----------------------------------
m
Bvhum Rham)1 4
jRSht  B)QRS5
S)t1 :hRRFLFDMCNRR:=w1qp S;
S)p1 :hRRFLFDMCNRR:=a )z
;S2
mSu)5aR
7SSjRR:H#MR0D8_FOoH;S
S7:4RRRHM#_08DHFoOS;
SR7.:MRHR8#0_oDFH
O;SdS7RH:RM0R#8F_Do;HO
7SScRR:H#MR0D8_FOoH;S
S7:6RRRHM#_08DHFoOS;
SR7n:MRHR8#0_oDFH
O;S(S7RH:RM0R#8F_Do;HO
7SSURR:H#MR0D8_FOoH;S
S7:gRRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SBSup:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SpwBiRR:H#MR0D8_FOoH;S
STRR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1)R4j:FRBlMbFCRM0H0#Rs;kC
--------------------7Qm Ypq---------------------------------
--
vBmu mhhQaRmp7 q
YRSht  B)QRR5RBa_1qBaQ_Y7pRH:RMo0CC:sR=2Rj;u
SmR)a5S
S7:QRRRQh#_08DHFoOS;
Sa17q:uRRRQh#_08DHFoOS;
Sa1 hRR:Q#hR0D8_FOoH;S
Sezqp RR:Q#hR0D8_FOoH;S
S7:mRRamzR8#0_oDFH
O;SwS7Rm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ m7pRqY:FRBlMbFCRM0H0#Rs;kC
--------------------vQ ---------------------------------
-
Bumvmhh a RQvSR
t  h)5QB
WSSQQh1Z: RRs#0HRMo:"=R1pvqp
";S1St)R h:FRLFNDCM=R:Rpwq1
 ;S1Sp)R h:FRLFNDCM=R:Rza) 2
S;u
SmR)a5S
S7RR:H#MR0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSvpRi:H#MR0D8_FOoH;S
SpRqt:kRF00R#8F_Do;HO
pSS Rq7:kRF00R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR :vRRlBFbCFMMH0R#sR0k
C;---------------------)--m-v--------------------------
-
Bumvmhh amR)vRR
RtRR )h Q5BRRR
SA_QaWaQ7]RR:HCM0oRCs:;=4SR
S)7 q_7vm RR:LRH0:'=Rj
';RRRRSpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRR
RRRRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
BSRpRi,Bm ,B) , a1 , W)RH:RM0R#8F_Do;HO
RRRRASRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
qSR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRm:vRRlBFbCFMMH0R#sR0k
C;-----------------------------m-)vRXg---------------------------------------------B

mmvuha hRv)mX
gRRRRRt  h)RQB5RR
RARRQWa_Q]7aRH:RMo0CC:sR=
g;RRRR)7 q_7vm RR:LRH0:j=''R;
RARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RRRRRRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
R
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoOR;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRv)mX:gRRlBFbCFMMH0R#sR0k
C;-----------------1--u---------------------------------------
m
Bvhum Rha1
uRRRRRt  h)RQB5R
SA_QaWaQ7]RR:HCM0oRCs:.=d;-R-RR4,.c,R,,RUR,4nR
d.S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SWa)Q m_v7: RR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRRaAY h_ q Ap_:jRR0LHRR:=';4'-j-''8:RHL#NDICRsCH0R:r(jL9RHR0;':4'RNCMLRDCI0sHC(Rr:Rj9L
H0RRRRRaAY h_ q Ap_:4RR0LHRR:=';4'-r-R4U6:9R
RRARRY_a  Ahqp. _RL:RH:0R=4R''-;-Rdr.:94n
RRRRYRAa  _hpqA R_d:HRL0=R:R''4;R--r:d4.
c9SpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"R
RRRRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
BSRpRi,Bm ,B) , a1 , W)RH:RM0R#8F_Do;HO
qSR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRRRSA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
S7:QRRRHM#_08DHFoOC_POs0F5Rd48MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV1:uRRlBFbCFMMH0R#sR0k
C;----------------------------1guX-------------------------------------
--
vBmu mhh1aRuRXg
RRRRht  B)QR
5RSQRAaQ_W7Ra]:MRH0CCos=R:gS;
Rq) 7m_v7: RR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
WSR) Qa_7vm RR:L_H0P0COF:sR=j"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRARRY_a  Ahqpj _RL:RH:0R=4R''-;-':j'R#8HNCLDRHIs0rCRU9:jR0LH;4R''C:RMDNLCsRIHR0CrjU:9HRL0R
RRARRY_a  Ahqp4 _RL:RH:0R=4R''-;-R(r4:
g9RRRRRaAY h_ q Ap_:.RR0LHRR:=';4'-r-R.4n:UR9
RRRRA Ya_q hA_p dRR:LRH0:'=R4-';-dRr6(:.9R
SA_pi1R p:HRL0C_POs0FRR:="jjj"S;
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRR
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoOS;
RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R;j2
RRRRASRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R
j2
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF1VRuRXg:FRBlMbFCRM0H0#Rs;kC
--------------------------------1--7-u--------------------------------------B

mmvuha hRu17RR
RR RthQ )BRR5
ASRQWa_Q]7a_:jRR0HMCsoCR4:=n-;R-,R4RR.,cU,R,nR4,.Rd
ASRQWa_Q]7a_:4RR0HMCsoCR4:=n-;R-,R4RR.,cU,R,nR4,.Rd
)SR _q7v m7RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8RC
RRRRA Ya_q hA_p jRR:LRH0:'=R4-';-''j:HR8#DNLCsRIHR0Crj(:9HRL0';R4R':CLMNDICRsCH0R:r(jL9RHR0
RRRRA Ya_q hA_p 4RR:LRH0:'=R4-';-4Rr69:U
RRRRYRAa  _hpqA R_.:HRL0=R:R''4;R--r:.d4
n9RRRRRaAY h_ q Ap_:dRR0LHRR:=';4'-r-Rd.4:cS9
RiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";ShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu17RB:RFFlbM0CMRRH#0Csk;-
---------------------------------1X7ug---------------------------------------
m
Bvhum Rha1X7ugRR
RtRR )h Q5BRRR
SA_QaWaQ7]R_j:MRH0CCos=R:4RU;-g-R,UR4,nRd
ASRQWa_Q]7a_:4RR0HMCsoCR4:=U-;R-,RgR,4UR
dnS R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SA Ya_q hA_p jRR:LRH0:'=R4-';-''j:HR8#DNLCsRIHR0CrjU:9HRL0';R4R':CLMNDICRsCH0R:rUjL9RHR0
RRRRA Ya_q hA_p 4RR:LRH0:'=R4
';RRRRRaAY h_ q Ap_:.RR0LHRR:=';4'
RRRRYRAa  _hpqA R_d:HRL0=R:R''4;R
SA_pi1R p:HRL0C_POs0FRR:="jjj"S;
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
RRRRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
BSRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  ,aAWq) , W)ARR:H#MR0D8_FOoH;R
Sq,7qqR7A:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;RRRRSpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7R1uRXg:FRBlMbFCRM0H0#Rs;kC
-----------------------------7u-------------------------------------
-
Bumvmhh auR7RR
RR RthQ )B
R5SASRQWa_Q]7a_:jRR0HMCsoCR4:=n
;RSASRQWa_Q]7a_:4RR0HMCsoCR4:=n
;RS)SR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)SR _q7v m74RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSWSR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CSWSR) Qa_7vm :4RR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRSYRAa  _hpqA __qjRR:LRH0:'=R4-';-''j:HR8#DNLCsRIHR0Cb0FsRrqR(9:jR0LH;4R''C:RMDNLCsRIHR0Crj(:9HRL0R
RRRRRRARRY_a  Ahqpq __:4RR0LHRR:=';4'-I-RsCH0RsbF0RRqr:46UR9
RRRRRRRRA Ya_q hA_p AR_j:HRL0=R:R''4;R--':j'R#8HNCLDRHIs0bCRFRs0A(Rr:Rj9L;H0R''4:MRCNCLDRHIs0rCR(9:jR0LH
RRRRRRRRYRAa  _hpqA __A4RR:LRH0:'=R4-';-sRIHR0Cb0FsRrAR4U6:9R
SRRRRSpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RSSQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
j"RRRR2R;
RuRRmR)a5S
SRq7m,A7mRF:Rk#0R0D8_FOoH_OPC05Fs486RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,42S;
SpRBiBq,p,iARqB ,AB , mBqB,m )A, a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRSRSRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuRR:BbFlFMMC0#RHRk0sC-;
-------------------------7--u-Xg-------------------------------------
-
Bumvmhh auR7X
gRRRRRt  h)RQB5SR
RaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUR
SA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4
)SR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
RQW)av _mj7 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
SWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RRRRYRAa  _hpqA __qjRR:LRH0:'=R4-';-''j:HR8#DNLCsRIHR0Cb0FsRrqRU9:jR0LH;4R''C:RMDNLCsRIHR0CrjU:9HRL0R
RRARRY_a  Ahqpq __:4RR0LHRR:=';4'-I-RsCH0RsbF0RRqr:4(gR9
RRRRA Ya_q hA_p AR_j:HRL0=R:R''4;'--jR':8NH#LRDCI0sHCFRbsA0RR:rUjL9RHR0;':4'RNCMLRDCI0sHCURr:Rj9L
H0RRRRRaAY h_ q Ap_4A_RL:RH:0R=4R''-;-RHIs0bCRFRs0A4Rr(9:g
RRRRASRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRR
RR;R2
RRRR)uma
R5SmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2O:=F_MP#_08DHFoOC_POs0F54j,U
2;SpRBiBq,p,iARqB ,AB , mBqB,m )A, a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
Rqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
7SRQ:qRRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2R;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RA7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR7X:gRRlBFbCFMMH0R#sR0k
C;--------------------------------)4qvn-14-------------------------B

mmvuha hRv)q44n1RR
RR RthQ )BRR5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jjRj"2R;
RuRRmR)a5S
S7:mRR0FkR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
SWR) :MRHR8#0_oDFH
O;S7SqjRR:H#MR0D8_FOoH;S
SqR74:MRHR8#0_oDFH
O;S7Sq.RR:H#MR0D8_FOoH;S
SqR7d:MRHR8#0_oDFH
O;SQS7RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n4RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41-.-------------------------
m
Bvhum Rha)4qvnR1.
RRRRht  B)QRQ5Rh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
"RRRRRRRRRRRRR2R;
RuRRmR)a5S
S7Rmj:kRF00R#8F_Do;HO
7SSm:4RR0FkR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
SWR) :MRHR8#0_oDFH
O;S7SqjRR:H#MR0D8_FOoH;S
SqR74:MRHR8#0_oDFH
O;S7Sq.RR:H#MR0D8_FOoH;S
SqR7d:MRHR8#0_oDFH
O;SQS7jRR:H#MR0D8_FOoH;S
S7RQ4:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRv)q4.n1RB:RFFlbM0CMRRH#0Csk;-
------------------------------q-)v14nc------------------------
--
vBmu mhh)aRqnv41
cRRRRRt  h)5QBRQQhaR_j:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
SRRRRQahQ_:4RR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RSRRQRRh_Qa.RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";RRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj
RRRRRRRRRRR2R;
RuRRmR)a5S
S7Rmj:kRF00R#8F_Do;HORS
S7Rm4:kRF00R#8F_Do;HO
7SSm:.RR0FkR8#0_oDFH
O;SmS7dRR:FRk0#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
Sjq7RH:RM0R#8F_Do;HO
qSS7:4RRRHM#_08DHFoOS;
S.q7RH:RM0R#8F_Do;HO
qSS7:dRRRHM#_08DHFoOS;
Sj7QRH:RM0R#8F_Do;HO
7SSQ:4RRRHM#_08DHFoOS;
S.7QRH:RM0R#8F_Do;HO
7SSQ:dRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnR1c:FRBlMbFCRM0H0#Rs;kC
--------------------------------v)q47n1u-4-------------------------

RRBumvmhh aqR)v14n7Ru4
RRRRht  B)Q5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj";R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S)SW RR:H#MR0D8_FOoH;S
SWjq7RH:RM0R#8F_Do;HO
WSSqR74:MRHR8#0_oDFH
O;SqSW7:.RRRHM#_08DHFoOS;
S7WqdRR:H#MR0D8_FOoH;S
S)jq7RH:RM0R#8F_Do;HO
)SSqR74:MRHR8#0_oDFH
O;SqS)7:.RRRHM#_08DHFoOS;
S7)qdRR:H#MR0D8_FOoH;S
S7:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu174RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41.7u-------------------------
-
Bumvmhh aqR)v14n7Ru.
RRRRht  B)QRQ5Rh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjjR"
RRRRRRRRR2RR;R
RRmRu)5aR
7SRm:jRR0FkR8#0_oDFH
O;SmR74RR:FRk0#_08DHFoOS;
RiBpRH:RM0R#8F_Do;HO
WSR): RRRHM#_08DHFoOS;
R7WqjRR:H#MR0D8_FOoH;R
SW4q7RH:RM0R#8F_Do;HO
WSRqR7.:MRHR8#0_oDFH
O;SqRW7:dRRRHM#_08DHFoOS;
R7)qjRR:H#MR0D8_FOoH;R
S)4q7RH:RM0R#8F_Do;HO
)SRqR7.:MRHR8#0_oDFH
O;SqR)7:dRRRHM#_08DHFoOS;
Rj7QRH:RM0R#8F_Do;HO
7SRQ:4RRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu17.RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41c7u-------------------------
-
Bumvmhh aqR)v14n7Ruc
RRRRht  B)QRQ5Rh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";RRRRRRRRRRRRRhRQQ.a_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R;
RRRRRRRRRRRRRQQhaR_d:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj
RRRRRRRRRRRR
2;RRRRuam)RS5
Sj7mRF:Rk#0R0D8_FOoH;S
S7Rm4:kRF00R#8F_Do;HO
7SSm:.RR0FkR8#0_oDFH
O;SmS7dRR:FRk0#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
S7WqjRR:H#MR0D8_FOoH;S
SW4q7RH:RM0R#8F_Do;HO
WSSqR7.:MRHR8#0_oDFH
O;SqSW7:dRRRHM#_08DHFoOS;
S7)qjRR:H#MR0D8_FOoH;S
S)4q7RH:RM0R#8F_Do;HO
)SSqR7.:MRHR8#0_oDFH
O;SqS)7:dRRRHM#_08DHFoOS;
Sj7QRH:RM0R#8F_Do;HO
7SSQ:4RRRHM#_08DHFoOS;
S.7QRH:RM0R#8F_Do;HO
7SSQ:dRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu17cRR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--mnv4-----------------------------B

mmvuha hRv)m4
nRRRRRt  h)RQB5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj";R2
RRRR)uma
R5R7SRmRR:FRk0#_08DHFoOS;
RRQj:MRHR8#0_oDFH
O;RRRRRRRRRRQ4:MRHR8#0_oDFH
O;S.RQRH:RM0R#8F_Do;HO
QSRdRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRmnv4RB:RFFlbM0CMRRH#0Csk;-
------------------A--z-wt-------------------------
-
Bumvmhh azRAw
tRRmRu)
a5RRRRS:mRR0FkR8#0_oDFH
O;RRRRS:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVAtzwRB:RFFlbM0CMRRH#0Csk;-
--------------A--z-w1-----------------
--
vBmu mhhAaRzRw1
RRRR)uma
R5RRRRRRRRR:mRR0FkR8#0_oDFH
O;RRRRRRRRR:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVA1zwRB:RFFlbM0CMRRH#0Csk;-
---------------------t-h7----------------
m
Bvhum RhatRh7
RRRR)uma
R5RRRRSRRt:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVhRt7RR:BbFlFMMC0#RHRk0sC-;
--------------------e-BB---------------------
--
vBmu mhheaRB
BRRRRRuam)RR5
RSRRR:eRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRBeBRB:RFFlbM0CMRRH#0Csk;-
-----------------m-1B-------------------------
--
vBmu mhhmaR1
BRRRRRuam)RS5
R1)  RaR:MRHR0R#8F_Do;HO
mSR1zBmaRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVmR1B:FRBlMbFCRM0H0#Rs;kC
----------------a-Kq-t------------------------------
--
vBmu mhhKaRaRqt
RRRR)uma
R5SaRK7RQR:kRF00R#8F_Do;HO
RRRRKSRaiBpRF:Rk#0R0D8_FOoH;R
SK1avRRR:FRk0#_08DHFoOR;
RRRRRRRRaR7mRRR:FRk0#_08DHFoOR;
RRRRRRRRaR7QRRR:HRMR#_08DHFoOR;
RRRRRRRRaiBpRRR:HRMR#_08DHFoOR;
RRRRRRRRaRv1RRR:HRMR#_08DHFoOR;
RRRRRRRRKma7RRR:HRMR#_08DHFoORRRRR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVKtaqRB:RFFlbM0CMRRH#0Csk;-
--------------Q--h-e------------------------------
--
vBmu mhhQaRh
eRRRRRuam)RR5
RSRRR:mRRamzR8#0_oDFH
O;RRRRSRRQ:hRQR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFReQhRB:RFFlbM0CMRRH#0Csk;-

----------------7-pp--------------------------------
vBmu mhh7aRpRp
RtRR )h Q
B5RRRRRRRR7_ppwBm) RR:HCM0oRCs:j=R;4--:FRVsROCD	FOR8NMR8OFCj;R:FRO8DC/FRO	oCCMsCN08sRVF7lRpDpRF
FbRRRRRRRRBQpihp1 R1:Rah)Qt=R:Rj"jj"j4;j--jjjj:#P#5V8CN0kD2j;jj:j4BQpihj;jj,4jjjj4j4,jj,jj4jjjjB:]phiQr~j9r
d9RRRRRRRR7_Qe1R p:HRL0=R:R''4;j--,sMFlRNDD	FOR8lFC4;R,#VN0FRDOl	RF
8CSRRRR7Bm q1BpRR:1Qa)h:tR=jR"j;j"-j-j44Rjj4Rj4jR4jjR444R4j4R44R
RRRRRRBR1q p_hRR:1Qa)h:tR=0R"s"kC-s-0kVC,NCD#
RRRR
2;RRRRuam)5R
RRRRRRBR]phiQRQ:Rh0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRBQpihh:QR8#0_oDFH=O:';j'
RRRRRRRRm1auQ:RM0R#8F_Do:HO=''j;R
RRRRRR R)1R a:MRQR8#0_oDFH=O:';j'
RRRRRRRR7zuhaBhpRR:Q#MR0D8_FOoH:j=''R;
RRRRRpRRmRBi:zRma0R#8F_Do;HO
RRRRRRRR 1auRR:mRza#_08DHFoOC_POs0F58(RF0IMF2Rj
RRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rpp:FRBlMbFCRM0H0#Rs;kC
-
--------------p--e_71QwAz---------------------------------B

mmvuha hR7pe1A_QzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7_zQAwRR:BbFlFMMC0#RHR""Q;-

----------------p1e7_zmAw--------------------------------
-
Bumvmhh aeRp7m1_A
zwRRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRR:QRRRQh#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRe_71mwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7pe1A_mz:wRRlBFbCFMMH0R#mR""
;
-----------------7pe1A_az-w------------------------------
--
vBmu mhhpaRe_71awAz
RRRR)umaR5
RRRRRmRRRm:Rz#aR0D8_FOoH;R
RRRRRRRRQ:hRQR8#0_oDFH
O;RRRRRRRRm: RRRQh#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRe_71awAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7pe1A_az:wRRlBFbCFMMH0R#mR""
;
-----------------7pe1m_QA-zw--------------------------------
m
Bvhum Rhap1e7_AQmzRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSQ:mRRmQhz#aR0D8_FOoH;R
RRSRRRRQR:hRQRRRR#_08DHFoOS;
RRRRRRm :hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRe_71QzmAwRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVeRp7Q1_mwAzRB:RFFlbM0CMRRH#"Rm,Q;m"
-
--------------p--e_71Atzw---------------------------------B

mmvuha hR7pe1z_AwRt
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp7A1_zRwt:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7_wAztRR:BbFlFMMC0#RHR""Q;-

----------------p1e7_wAz1--------------------------------
-
Bumvmhh aeRp7A1_z
w1RRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRR:QRRRQh#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRe_71A1zwRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7pe1z_Aw:1RRlBFbCFMMH0R#QR""
;
-----------------7pe1_.6QwAz---------------------------------B

mmvuha hR7pe1_.6QwAz
RRRR)umaR5
RRRRRmRRRm:Rz#aR0D8_FOoH;R
RRRRRRRRQ:hRQR8#0_oDFH
O;RRRRRRRRQ:ARRRQh#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRe.716A_Qz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFpVRe.716A_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------7pe1_ddQwAz---------------------------------B

mmvuha hR7pe1_ddQwAz
RRRR)umaR5
RRRRRmRRRm:Rz#aR0D8_FOoH;R
RRRRRRRRQ:hRQR8#0_oDFH
O;RRRRRRRRQ:ARRRQh#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRed71dA_Qz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFpVRed71dA_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------7pe1_.6mwAz---------------------------------B

mmvuha hR7pe1_.6mwAz
RRRR)umaR5
RRRRRmRRRm:Rz#aR0D8_FOoH;R
RRRRRRARmRm:Rz#aR0D8_FOoH;R
RRRRRRRRQ:hRQR8#0_oDFHRO
RRRRR2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVp1e7.m6_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7.m6_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------e-p7d1d_zmAw--------------------------------
-
Bumvmhh aeRp7d1d_zmAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRmRRARR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFR7pe1_ddmwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7pe1_ddmwAzRB:RFFlbM0CMRRH#"Rm,m;A"R
RR
----------------e-p761._zaAw--------------------------------
-
Bumvmhh aeRp761._zaAwR
RRmRu)5aR
RRRRmSRRRR:mRzaR0R#8F_Do;HO
RRRRmSRARR:mRza#_08DHFoOR;
RRRRSRRQRQ:RhRRRR8#0_oDFH
O;SRRRR RmRQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVp1e7.a6_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7.a6_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------e-p7d1d_zaAw--------------------------------
-
Bumvmhh aeRp7d1d_zaAwR
RRmRu)5aR
RRRRmSRRRR:mRzaR0R#8F_Do;HO
RRRRmSRARR:mRza#_08DHFoOR;
RRRRSRRQRQ:RhRRRR8#0_oDFH
O;SRRRR RmRQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVp1e7dad_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7dad_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------e-p761._AQmz-w------------------------------
--
vBmu mhhpaRe.716m_QA
zwRRRRuam)RR5
RSRRRRmR:zRmaRRR#_08DHFoOR;
RSRRRAQmRQ:RhamzR8#0_oDFH
O;RRRRRRRRRRQm:hRQmRza#_08DHFoOR;
RRRRSRRQRQ:RhRRRR8#0_oDFH
O;SRRRR RmRQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVp1e7.Q6_mwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFR7pe1_.6QzmAwRR:BbFlFMMC0#RHR,"mR,QmRAQm"
;
-----------------7pe1_ddQzmAw--------------------------------
-
Bumvmhh aeRp7d1d_AQmzRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSQRmA:hRQmRza#_08DHFoOR;
RRRRRRRRQ:mRRmQhz#aR0D8_FOoH;R
RRSRRRRQR:hRQRRRR#_08DHFoOS;
RRRRRRm :hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFpVRed71dm_QARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVp1e7dQd_mwAzRB:RFFlbM0CMRRH#"Rm,QRm,Q"mA;-

----------------p1e7.A6_z-wt--------------------------------
m
Bvhum Rhap1e7.A6_z
wtRRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp761._wAztRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVeRp761._wAztRR:BbFlFMMC0#RHR,"QR"QA;-

----------------p1e7dAd_z-wt--------------------------------
m
Bvhum Rhap1e7dAd_z
wtRRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp7d1d_wAztRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVeRp7d1d_wAztRR:BbFlFMMC0#RHR,"QR"QA;-

----------------p1e7.A6_z-w1--------------------------------
m
Bvhum Rhap1e7.A6_z
w1RRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp761._wAz1RR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVeRp761._wAz1RR:BbFlFMMC0#RHR,"QR"QA;-

----------------p1e7dAd_z-w1--------------------------------
m
Bvhum Rhap1e7dAd_z
w1RRRRuam)5R
RRRRRRRRm:zRma0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVeRp7d1d_wAz1RR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVeRp7d1d_wAz1RR:BbFlFMMC0#RHR,"QR"QA;RRRR-

-------------------------v--z4paUUX47---------------------------------------
vBmu mhhvaRz4paUUX47S
SoCCMs5HO
RSSRQRRh)q_ :tRRHRL0=R:R''j;-R-RjR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
RSSRQRRh)A_ :tRRHRL0=R:R''j;S
SRRRRm_za)R t:LRRH:0R=jR''S;
SRRRRuuQ  _)tRR:R0LHRR:=';j'
RSSRqRR1hQt__Qh)R t:LRRH:0R=jR''S;
SRRRRQq1tuh_Q_u )R t:LRRH:0R=jR''S;
SRRRRQA1tQh_h _)tRR:R0LHRR:=';j'
RSSRARR1hQt_uuQ  _)tRR:R0LHRR:=';j'
RSSRvRRz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"-R-Rh1YBq,R1BYh
RSRR;R2
RRRRRRR
RRRRRRRR)umaS5
S7SvQ:qRRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SRRRRQv7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SRRRRqt1QhA,R1hQtRH:RM0R#8F_Do;HO
RSSRBRR RR:H#MR0D8_FOoH;S
SRRRRBRpi:MRHR8#0_oDFH
O;SRSRR R)1R a:MRHR8#0_oDFH
O;SRSRRmRvz:aRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;SRSRR1RvQRth:kRF00R#8F_Do
HOS;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazp44UXU:7RRlBFbCFMMH0R#sR0k
C;
----------------------------pvzaggX7---------------------------------------
m
Bvhum Rhavazpg7Xg
RRRRMoCCOsH5S
SRRRRQ_hq)R t:LRRH:0R=jR''-;R-'RRjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SRRRRQ_hA)R t:LRRH:0R=jR''S;
SRRRRamz_t) RR:RLRH0:'=Rj
';SRSRRQRuu) _ :tRRHRL0=R:R''j;S
SRRRRqt1Qhh_Q_t) RR:RLRH0:'=Rj
';SRSRR1RqQ_thu Qu_t) RR:RLRH0:'=Rj
';SRSRR1RAQ_thQ)h_ :tRRHRL0=R:R''j;S
SRRRRAt1QhQ_uu) _ :tRRHRL0=R:R''j;S
SRRRRvazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YBR
SR2RR;R
RRRRRRSR
b0FsRS5
SRRRRQv7qRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
RSSRvRR7RQA:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SRRRRQq1tRh,At1QhRR:H#MR0D8_FOoH;S
SRRRRB: RRRHM#_08DHFoOS;
SRRRRiBpRH:RM0R#8F_Do;HO
RSSR)RR a1 RH:RM0R#8F_Do;HO
RSSRvRRmRza:kRF00R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
RSSRvRR1hQtRF:Rk#0R0D8_FOoH
RSRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpg7XgRB:RFFlbM0CMRRH#0Csk;-

-------------------------v--z4paUUX41------------------------------------B-
mmvuha hRpvzaX4U4
U1SCSoMHCsOS5
SqQh_t) RR:RLRH0:'=RjR';-R-R':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SAQh_t) RR:RLRH0:'=Rj
';SzSma _)tRR:R0LHRR:=';j'
uSSQ_u )R t:LRRH:0R=jR''S;
SQq1tQh_h _)tRR:R0LHRR:=';j'
qSS1hQt_uuQ  _)tRR:R0LHRR:=';j'
ASS1hQt__Qh)R t:LRRH:0R=jR''S;
SQA1tuh_Q_u )R t:LRRH:0R=jR''R;
RRRRR1RR]aQw_amz_t) RL:RH:0R=jR''S;
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2R;
R
RRSsbF0
R5S7SvQ1q,7RQq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;S7SvQ1A,7RQA:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;S1SqQ,thRQA1t:hRRRHM#_08DHFoOR;
RRRRRqRR1, pR A1pRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
vSSmRza:kRF00R#8F_Do_HOP0COFds56FR8IFM0R;j2
RRRRRRRRm17q7,1m:ARR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;S1SvQRth:kRF00R#8F_Do
HOS
2; Rh7Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz4paUUX41RR:BbFlFMMC0#RHRk0sC
;
----------------------------vazpg1Xg-------------------------------------
--
vBmu mhhvaRzgpaX
g1RRRRoCCMs5HO
QSSh)q_ :tRRHRL0=R:R''j;-R-RjR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
QSSh)A_ :tRRHRL0=R:R''j;S
Sm_za)R t:LRRH:0R=jR''S;
SuuQ  _)tRR:R0LHRR:=';j'
qSS1hQt__Qh)R t:LRRH:0R=jR''S;
SQq1tuh_Q_u )R t:LRRH:0R=jR''S;
SQA1tQh_h _)tRR:R0LHRR:=';j'
ASS1hQt_uuQ  _)tRR:R0LHRR:=';j'
RRRRRRRRQ1]wma_z)a_ :tRRHRL0=R:R''j;SR
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5S7SvQ1q,7RQq:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SQv7A7,1Q:ARRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
Sqt1QhA,R1hQtRH:RM0R#8F_Do;HO
RRRRRRRR q1p1,A :pRRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SvamzRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj;R
RRRRRR7R1m1q,7RmA:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;S1SvQRth:kRF00R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzgpaXRg1:FRBlMbFCRM0H0#Rs;kC
-
--------------------------z-vpnadX74U-------------------------------------
--Bumvmhh azRvpnadX74U
CSoMHCsOS5
SRRRRqQh_t) RR:RLRH0:'=RjR';-R-R':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SRRRRAQh_t) RR:RLRH0:'=Rj
';SRSRRzRma _)tRR:R0LHRR:=';j'
RSSRuRRQ_u )R t:LRRH:0R=jR''S;
SRRRRQq1tQh_h _)tRR:R0LHRR:=';j'
RSSRqRR1hQt_uuQ  _)tRR:R0LHRR:=';j'
RSSRARR1hQt__Qh)R t:LRRH:0R=jR''S;
SRRRRQA1tuh_Q_u )R t:LRRH:0R=jR''S;
SRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
RRRR2R;
RRRRR
RRSsbF0
R5S7SvQ:qRRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
SQv7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
Sqt1QhA,R1hQtRH:RM0R#8F_Do;HO
BSS RR:H#MR0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;RRRRRRRRvt1QhRR:FRk0#_08DHFoOS;
SzvmaRR:FRk0#_08DHFoOC_POs0F5R6d8MFI0jFR22
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvzaXdn4RU7:FRBlMbFCRM0H0#Rs;kC
-
--------------------------z-vpnadX7dn-------------------------------------
--Bumvmhh azRvpnadX7dn
CSoMHCsOS5
SRRRRqQh_t) RR:RLRH0:'=RjR';-R-R':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SRRRRAQh_t) RR:RLRH0:'=Rj
';SRSRRzRma _)tRR:R0LHRR:=';j'
RSSRuRRQ_u )R t:LRRH:0R=jR''S;
SRRRRQq1tQh_h _)tRR:R0LHRR:=';j'
RSSRqRR1hQt_uuQ  _)tRR:R0LHRR:=';j'
RSSRARR1hQt__Qh)R t:LRRH:0R=jR''S;
SRRRRQA1tuh_Q_u )R t:LRRH:0R=jR''S;
SRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
RRRR2S;

FSbs50R
vSS7RQq:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;S7SvQ:ARRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
SQq1tRh,At1QhRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
RRRRRRRR1vQt:hRR0FkR8#0_oDFH
O;SmSvz:aRR0FkR8#0_oDFHPO_CFO0s45(RI8FMR0FjS2
2 ;
hB7Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvpnadX7dnRB:RFFlbM0CMRRH#0Csk;R
RR-R
-------------------------v--zqpa7U74X74U-------------------------------------
--Bumvmhh azRvp7aq7X4U4
U7SMoCCOsH5S
SQjhq_t) RL:RH:0R=jR''-;-R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CShSQA)j_ :tRR0LHRR:=';j'RS
SQ4hq_t) RL:RH:0R=jR''S;
SAQh4 _)tRR:LRH0:'=Rj
';SzSma _)tRR:LRH0:'=Rj
';SQSuu_ j)R t:HRL0=R:R''j;S
Su Qu4 _)tRR:LRH0:'=Rj
';S1SqQjth__Qh)R t:HRL0=R:R''j;S
SAt1QhQj_h _)tRR:LRH0:'=Rj
';S1SqQ4th__Qh)R t:HRL0=R:R''j;S
SAt1QhQ4_h _)tRR:LRH0:'=Rj
';S1SqQjth_uuQ  _)tRR:LRH0:'=Rj
';S1SAQjth_uuQ  _)tRR:LRH0:'=Rj
';S1SqQ4th_uuQ  _)tRR:LRH0:'=Rj
';S1SAQ4th_uuQ  _)tRR:LRH0:'=Rj
';S7Sq7A1z_t) jRR:LRH0:'=Rj
';S7Sq7A1z_t) 4RR:LRH0:'=Rj
';SzSvp)a_ a1 _7vm RR:#H0sM:oR=1R"Y"hBRR--1BYh,1RqY
hBS
2;
FSbs50R
vSS7jQq,Qv7q:4RRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SQv7Avj,74QARH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
RRRRRRRRQq1tRh,At1QhRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RRRRRRRR7q71RzA:MRHR8#0_oDFH
O;S SBRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SzvmaRR:FRk0#_08DHFoOC_POs0F5Rdn8MFI0jFR22
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvza7q744UXU:7RRlBFbCFMMH0R#sR0k
C;
----------------------------pvza7q7g7Xg-------------------------------------
--Bumvmhh azRvp7aq7ggX7o
SCsMCH
O5ShSQq)j_ :tRR0LHRR:=';j'-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SQjhA_t) RL:RH:0R=jR''
;RShSQq)4_ :tRR0LHRR:=';j'
QSSh_A4)R t:HRL0=R:R''j;S
Sm_za)R t:HRL0=R:R''j;S
Su Quj _)tRR:LRH0:'=Rj
';SQSuu_ 4)R t:HRL0=R:R''j;S
Sqt1QhQj_h _)tRR:LRH0:'=Rj
';S1SAQjth__Qh)R t:HRL0=R:R''j;S
Sqt1QhQ4_h _)tRR:LRH0:'=Rj
';S1SAQ4th__Qh)R t:HRL0=R:R''j;S
Sqt1Qhuj_Q_u )R t:HRL0=R:R''j;S
SAt1Qhuj_Q_u )R t:HRL0=R:R''j;S
Sqt1Qhu4_Q_u )R t:HRL0=R:R''j;S
SAt1Qhu4_Q_u )R t:HRL0=R:R''j;S
Sq177z)A_ Rtj:HRL0=R:R''j;S
Sq177z)A_ Rt4:HRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
SQv7qvj,74QqRH:RM0R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;S7SvQ,AjvA7Q4RR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
RRRRRRRRQq1tRh,At1QhRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RRRRRRRR7q71RzA:MRHR8#0_oDFH
O;S SBRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SzvmaRR:FRk0#_08DHFoOC_POs0F5R4U8MFI0jFR22
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvza7q7g7XgRB:RFFlbM0CMRRH#0Csk;-

-------------------------v--zqpa7z71vX4U4-U7-------------------------------------B-
mmvuha hRpvza7q714zvUUX47o
SCsMCH
O5ShSQq)j_ :tRR0LHRR:=';j'RR--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SAQhj _)tRR:LRH0:'=RjR';
QSSh_q4)R t:HRL0=R:R''j;SR
SAQh4 _)tRR:LRH0:'=RjR';
RRRRRRRRqQh. _)tRR:LRH0:'=RjR';
QSSh_A.)R t:HRL0=R:R''j;RR
RRRRRQRRh_qd)R t:HRL0=R:R''j;SR
SAQhd _)tRR:LRH0:'=RjR';
RRRRRRRRamz_t) RL:RH:0R=jR''S;
SuuQ )j_ :tRR0LHRR:=';j'
uSSQ4u _t) RL:RH:0R=jR''S;
SuuQ )._ :tRR0LHRR:=';j'
uSSQdu _t) RL:RH:0R=jR''S;
SQq1t_hjQ)h_ :tRR0LHRR:=';j'
qSS1hQtjQ_uu) _ :tRR0LHRR:=';j'
ASS1hQtjh_Q_t) RL:RH:0R=jR''S;
SQA1t_hju Qu_t) RL:RH:0R=jR''S;
SQq1t_h4Q)h_ :tRR0LHRR:=';j'
qSS1hQt4Q_uu) _ :tRR0LHRR:=';j'
ASS1hQt4h_Q_t) RL:RH:0R=jR''S;
SQA1t_h4u Qu_t) RL:RH:0R=jR''S;
SQq1t_h.Q)h_ :tRR0LHRR:=';j'
qSS1hQt.Q_uu) _ :tRR0LHRR:=';j'
ASS1hQt.h_Q_t) RL:RH:0R=jR''S;
SQA1t_h.u Qu_t) RL:RH:0R=jR''S;
SQq1t_hdQ)h_ :tRR0LHRR:=';j'
qSS1hQtdQ_uu) _ :tRR0LHRR:=';j'
ASS1hQtdh_Q_t) RL:RH:0R=jR''S;
SQA1t_hdu Qu_t) RL:RH:0R=jR''R;
RRRRRqRR7z71A)j_ Rtj:HRL0=R:R''j;R
RRRRRR7Rq7A1zj _)t:4RR0LHRR:=';j'
RRRRRRRR7q714zA_t) jRR:LRH0:'=Rj
';RRRRRRRRq177z_A4)4 tRL:RH:0R=jR''S;
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5S7SvQ,qjvq7Q47,vQ,q.vq7QdRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SvA7Qj7,vQ,A4vA7Q.7,vQRAd:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;RRRRRRRRqt1QhA,R1hQtRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRq177z:ARRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
vSSmRza:kRF00R#8F_Do_HOP0COFds5(FR8IFM0R
j2S
2; Rh7Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzqpa7z71vX4U4RU7:FRBlMbFCRM0H0#Rs;kC
-
--------------------------z-vp7aq7v1zg7Xg-------------------------------------
--Bumvmhh azRvp7aq7v1zg7Xg
CSoMHCsOS5
SqQhj _)tRR:LRH0:'=RjR';-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SQjhA_t) RL:RH:0R=jR''
;RShSQq)4_ :tRR0LHRR:=';j'RS
SQ4hA_t) RL:RH:0R=jR''
;RRRRRRRRRQ.hq_t) RL:RH:0R=jR''
;RShSQA)._ :tRR0LHRR:=';j'RR
RRRRRRhRQq)d_ :tRR0LHRR:=';j'RS
SQdhA_t) RL:RH:0R=jR''
;RRRRRRRRRm_za)R t:HRL0=R:R''j;S
Su Quj _)tRR:LRH0:'=Rj
';SQSuu_ 4)R t:HRL0=R:R''j;S
Su Qu. _)tRR:LRH0:'=Rj
';SQSuu_ d)R t:HRL0=R:R''j;S
Sqt1QhQj_h _)tRR:LRH0:'=Rj
';S1SqQjth_uuQ  _)tRR:LRH0:'=Rj
';S1SAQjth__Qh)R t:HRL0=R:R''j;S
SAt1Qhuj_Q_u )R t:HRL0=R:R''j;S
Sqt1QhQ4_h _)tRR:LRH0:'=Rj
';S1SqQ4th_uuQ  _)tRR:LRH0:'=Rj
';S1SAQ4th__Qh)R t:HRL0=R:R''j;S
SAt1Qhu4_Q_u )R t:HRL0=R:R''j;S
Sqt1QhQ._h _)tRR:LRH0:'=Rj
';S1SqQ.th_uuQ  _)tRR:LRH0:'=Rj
';S1SAQ.th__Qh)R t:HRL0=R:R''j;S
SAt1Qhu._Q_u )R t:HRL0=R:R''j;S
Sqt1QhQd_h _)tRR:LRH0:'=Rj
';S1SqQdth_uuQ  _)tRR:LRH0:'=Rj
';S1SAQdth__Qh)R t:HRL0=R:R''j;S
SAt1Qhud_Q_u )R t:HRL0=R:R''j;R
RRRRRR7Rq7A1zj _)t:jRR0LHRR:=';j'
RRRRRRRR7q71jzA_t) 4RR:LRH0:'=Rj
';RRRRRRRRq177z_A4)j tRL:RH:0R=jR''R;
RRRRRqRR7z71A)4_ Rt4:HRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
SQv7qvj,74Qq,Qv7qv.,7dQqRH:RM0R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;S7SvQ,AjvA7Q47,vQ,A.vA7QdRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
RRRRRRRRQq1tRh,At1QhRR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRR7q71RzA:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SvamzRF:Rk#0R0D8_FOoH_OPC05Fs48gRF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpq177zXvgg:7RRlBFbCFMMH0R#sR0k
C;
----------------------------Bvq44UXU-7--------------------------------------m
Bvhum Rhav4qBUUX47o
SCsMCH
O5ShSQq _)tRR:LRH0:'=Rj-';-jR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
QSSh)A_ :tRR0LHRR:=';j'RS
Sp_7Q)_ tBRpi:HRL0=R:R''j;SR
S7q71_zA)j tRL:RH:0R=jR''
;RRRRRRRRRq177z)A_ Rt4:HRL0=R:R''j;RR
RRRRRqRRBmBpq)7_ Rtj:HRL0=R:R''j;R
RRRRRRBRqBqpm7 _)t:4RR0LHRR:=';j'
uSSQ_u )R t:HRL0=R:R''j;S
Sqt1Qhh_Q_t) RL:RH:0R=jR''S;
SQA1tQh_h _)tRR:LRH0:'=Rj
';S1SqQ_thu Qu_t) RL:RH:0R=jR''S;
SQA1tuh_Q_u )R t:HRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
SQv7qRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SvA7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
RRRRRRRRQq1tRh,At1QhRR:H#MR0D8_FOoH;R
RRRRRR7Rq7A1z,BRqBqpm7RR:H#MR0D8_FOoH;R
RRRRRR7RpQRR:H#MR0D8_FOoH_OPC05Fs68dRF0IMF2Rj;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
vSSmRza:kRF00R#8F_Do_HOP0COF6s5dFR8IFM0R;j2
RRRRRRRR me)mwpWRR:FRk0#_08DHFoO2
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRBvq44UXU:7RRlBFbCFMMH0R#sR0k
C;
----------------------------Bvqg7Xg-------------------------------------
--Bumvmhh aqRvBggX7o
SCsMCH
O5ShSQq _)tRR:LRH0:'=Rj-';-jR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
QSSh)A_ :tRR0LHRR:=';j'RS
Sp_7Q)_ tBRpi:HRL0=R:R''j;SR
S7q71_zA)j tRL:RH:0R=jR''
;RRRRRRRRRq177z)A_ Rt4:HRL0=R:R''j;RR
RRRRRqRRBmBpq)7_ Rtj:HRL0=R:R''j;R
RRRRRRBRqBqpm7 _)t:4RR0LHRR:=';j'
uSSQ_u )R t:HRL0=R:R''j;S
Sqt1Qhh_Q_t) RL:RH:0R=jR''S;
SQA1tQh_h _)tRR:LRH0:'=Rj
';S1SqQ_thu Qu_t) RL:RH:0R=jR''S;
SQA1tuh_Q_u )R t:HRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
SQv7qRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
vSS7RQA:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2R;
RRRRRqRR1hQt,1RAQRth:MRHR8#0_oDFH
O;RRRRRRRRq177zRA,qpBBmRq7:MRHR8#0_oDFH
O;RRRRRRRRpR7Q:MRHR8#0_oDFHPO_CFO0sn5.RI8FMR0Fj
2;S SBRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SzvmaRR:FRk0#_08DHFoOC_POs0F5R.n8MFI0jFR2R;
RRRRRmRRew )pRmW:kRF00R#8F_Do
HOS
2; Rh7Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRqXBgg:7RRlBFbCFMMH0R#sR0k
C;
----------------------------7uq7-4U-------------------------------------B-
mmvuha hR7uq7
4USMoCCOsH5S
SQ_hq)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SAQh_t) RL:RH:0R=jR''
;RShSQB _)tRR:LRH0:'=Rj
';S7Sq7A1z_t) RL:RH:0R=jR''R;
RRRRRuRRq_77)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-YR1hqB,1BYh
1SS]aQw_amz_t) RL:RH:0R=jR''R;
RRRRRqRR_1B_ :pRR0LHRR:=';j'RR--q
,BRRRRRRRRAp1 _7vm RR:L_H0P0COF:sR=4R"4R";-"-R4:4"RH#EVR0,""jj:NRbsDNDCHDRM0bkRQu7A",Rj:4"RqQh_t) 3R
RRRRRRARw__QhvRzX:HRL0=R:R''j;-R-R''j:ER#H,V0R''4:hRQq _)tR;
RRRRRQRRhvq_z:XRR0LHRR:='Rj'-'-R4R':#CCDOu0R7RQq8CHsO$0D;jR''Q:Rh)q_ 
t3S
2;
FSbs
05S7SuQ:qRRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SQu7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SuB7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
qSS1, pR7q71RzA:MRHR8#0_oDFH
O;S SB,iBp,1)  :aRRRHM#_08DHFoOS;
SQ17qq,u7Q71RH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
1SS7,mqu7q71:mRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SmSuz:aRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0FjS2
2 ;
hB7Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqRu7U74RB:RFFlbM0CMRRH#0Csk;-

-------------------------u--qg77-------------------------------------
--Bumvmhh aqRu7
7gSMoCCOsH5S
SQ_hq)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SAQh_t) RL:RH:0R=jR''
;RShSQB _)tRR:LRH0:'=Rj
';S7Sq7A1z_t) RL:RH:0R=jR''R;
RRRRRuRRq_77)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-YR1hqB,1BYh
1SS]aQw_amz_t) RL:RH:0R=jR''R;
RRRRRqRR_1B_ :pRR0LHRR:=';j'RR--q
,BRRRRRRRRAp1 _7vm RR:L_H0P0COF:sR=4R"4R";-"-R4:4"RH#EVR0,""jj:NRbsDNDCHDRM0bkRQu7A",Rj:4"RqQh_t) 3R
RRRRRRARw__QhvRzX:HRL0=R:R''j;-R-R''j:ER#H,V0R''4:hRQq _)tR;
RRRRRQRRhvq_z:XRR0LHRR:='Rj'-'-R4R':#CCDOu0R7RQq8CHsO$0D;jR''Q:Rh)q_ 
t3S
2;
FSbs
05S7SuQ:qRRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
SuA7QRH:RM0R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;S7SuQ:BRRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
Sqp1 ,7Rq7A1zRH:RM0R#8F_Do;HO
BSS p,Bi ,)1R a:MRHR8#0_oDFH
O;S7S1Quq,q177QRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
1SS7,mqu7q71:mRR0FkR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SzumaRR:FRk0#_08DHFoOC_POs0F58URF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVu7q7gRR:BbFlFMMC0#RHRk0sC
;
----------------------------q6pzc---------------------------------------
vBmu mhhqaRpcz6
CSoMHCsOS5
RRRRQ_hB)R t:HRL0=R:R''j;-R-':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
RRRRq1pz )p_ Rtj:HRL0=R:R''j;R
SRqRRp z1p _)t:4RR0LHRR:=';j'
RSRRpRqz7vm  _)t:jRR0LHRR:=';j'
RSRRpRqz7vm  _)t:4RR0LHRR:=';j'
RSRRzRma _)tRR:LRH0:'=Rj
';SRRRR_wA)R t:HRL0=R:R''j;R
SRvRRB)_1Bm_v7: RR0LHRR:=';j'RR--':j'RD#CCRO0vQB_h;QaR''4:D#CCRO0Q
hBSRRRR1vqi)_1Bm_v7: RR0LHRR:=';j'RR--':j'RD#CCRO0viq1_QQha';R4#':CODC0hRQBR
SRvRRqZ1imh_QQ:aRR0LH_OPC0RFs:X=R"jjjjjjjjjjjj"jj;R
SRvRRBh_QQ:aRR0LH_OPC0RFs:X=R"jjjjjjjjjjjj"jj;R
SRvRRq_1iQahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjj
";SRRRR7)h_QQhaRR:L_H0P0COF:sR="RXjjjjjjjjjjjjj;j"
RSRRpRqz _)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRvazpgm_v7: RR0LHRR:='Rj'-j-''l:Rk4D0UFRl8RC;':4'RDlk0lgRF
8CRRRR2R;
RbRRFRs05R
SRQRRh:qRRRHM#_08DHFoOC_POs0FR65dRI8FMR0Fj
2;SRRRRAQhRH:RM0R#8F_Do_HOP0COF5sRd86RF0IMF2Rj;R
SRwRRARR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRB: RRRHM#_08DHFoOS;
RRRRBRpi:MRHR8#0_oDFH
O;SRRRR1)  :aRRRHM#_08DHFoOS;
RRRRqt1Qh1,AQ,thBQQ1t:hRRRHM#_08DHFoOS;
RRRRQRhB:MRHR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
RSRR7RvjRR:H#MR0D8_FOoH_OPC0RFs5Rd68MFI0jFR2S;
RRRRvR74:MRHR8#0_oDFHPO_CFO0sdR56FR8IFM0R;j2
RSRRQRBhRR:H#MR0D8_FOoH_OPC0RFs5R6c8MFI0jFR2S;
RRRRq1pz :pRRRHM#_08DHFoOC_POs0F58nRF0IMF2Rj;R
RRRRRRpRqz7vm RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
RSRRmRBz:aRR0FkR8#0_oDFHPO_CFO0s6R5cFR8IFM0R;j2
RSRRARwB:mRR0FkR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
RSRRvRBuvZ,BZvu,vvBuvm,7uBv,hv7BRvu:kRF00R#8F_Do;HO
RSRReRm z),h)7 RF:Rk#0R0D8_FOoH;R
SRBRRmt1QhRR:FRk0#_08DHFoOR
RR;R2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVq6pzcRR:BbFlFMMC0#RHRk0sC
;
----------------------------q6pzc-]--------------------------------------m
Bvhum Rhaq6pzcS]
oCCMs5HO
RSRRhRQB _)tRR:LRH0:'=RjR';-j-''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
RSRRpRqzp1 _t) jRR:LRH0:'=Rj
';SRRRRzqp1_ p)4 tRL:RH:0R=jR''S;
RRRRqvpzm_7 )j tRL:RH:0R=jR''S;
RRRRqvpzm_7 )4 tRL:RH:0R=jR''S;
RRRRm_za)R t:HRL0=R:R''j;R
SRwRRA _)tRR:LRH0:'=Rj
';SRRRR_vB1_)Bv m7RL:RH:0R=jR''-;R-jR''#:RCODC0BRv_QQha';R4#':CODC0hRQBR
SRvRRq_1i1_)Bv m7RL:RH:0R=jR''-;R-jR''#:RCODC0qRv1Qi_h;QaR''4:D#CCRO0Q
hBSRRRR1vqi_ZmQahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjj
";SRRRR_vBQahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjj
";SRRRR1vqih_QQ:aRR0LH_OPC0RFs:X=R"jjjjjjjjjjjj"jj;R
SR)RRhQ7_hRQa:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjj"S;
RRRRq_pz)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRzRvp_agv m7RL:RH:0R=jR''-R-':j'RDlk0R4UlCF8;4R''l:RkgD0R8lFCR
RR;R2
RRRRsbF0
R5SRRRRqQhRH:RM0R#8F_Do_HOP0COF5sRd86RF0IMF2Rj;R
SRQRRh:ARRRHM#_08DHFoOC_POs0FR65dRI8FMR0Fj
2;SRRRRRwA:MRHR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
RSRR RBRH:RM0R#8F_Do;HO
RSRRpRBiRR:H#MR0D8_FOoH;R
SR)RR a1 RH:RM0R#8F_Do;HO
RSRR1RqQ,thAt1QhQ,B1hQtRH:RM0R#8F_Do;HO
RSRRhRQBRR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRvR7j:MRHR8#0_oDFHPO_CFO0sdR56FR8IFM0R;j2
RSRR7Rv4RR:H#MR0D8_FOoH_OPC0RFs5Rd68MFI0jFR2S;
RRRRBRQh:MRHR8#0_oDFHPO_CFO0s6R5cFR8IFM0R;j2
RSRRpRqzp1 RH:RM0R#8F_Do_HOP0COFns5RI8FMR0Fj
2;RRRRRRRRqvpzmR7 :MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
RRRR7amzRF:Rk#0R0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRBamzRF:Rk#0R0D8_FOoH_OPC0RFs5R6c8MFI0jFR2S;
RRRRwmABRF:Rk#0R0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRBZvu,vvBuvZ,Bmvu,Bv7vvu,7vhBuRR:FRk0#_08DHFoOS;
RRRRm)e ,7zh :)RR0FkR8#0_oDFH
O;SRRRR1BmQRth:kRF00R#8F_Do
HORRRR2 ;
hB7Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRqz]6cRB:RFFlbM0CMRRH#0Csk;R
RRRRRRRRRR-
------------------------------p-up------------------------
--Bumvmhh apRupR
RR RthQ )BR5
RRRRRRRRRRRRwiBpQ:hRR)1aQRht:"=R43jjjR";-s-VCCJkMRO$F0VREOCRDM	H5
v2RRRRRRRRRRRRRh7Y__Qh1R p:aR1)tQhRR:="DVN#;C"-s-0kQC:hp1 ;NRVD:#CR_Qh1
 pRRRRRRRRRRRRR_Qh1R p:MRH0CCos=R:R-6;-Bj:phiQr,694p:BirQhc.9,:iBpQdhr9:,dBQpih9r.,Bc:phiQr,496p:BirQhj89,CkVND
0RRRRRRRRRRRRRRh7Y_QQ7e _1pRR:1Qa)h:tR=VR"NCD#"-;-0Csk:1Q7 Rp;V#NDC7:QQ1e_ Rp
RRRRRRRRRRRRQe7Q_p1 RH:RMo0CC:sR=;Rj-M-QbRk08HHP8RCsQe7Q,:Rj4:,4.333nnd:cR3R4c~n
RRRRRRRRRRRRYR7hA_w7_Qe1R p:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRARw7_Qe1R p:MRH0CCos=R:R-j;-CwC8OLN	HR8PCH8sARw7,QeR:Rj4:,4.333nnd:c43R~
ncRRRRRRRRRRRRRQm7e _1pRR:HCM0oRCs:U=R;.--/Uc///4ndc./Uc/n//Ujg4n/44./.RU
RRRRRRRRRRRRuq17_p1 R1:Rah)Qt=R:Rj"jj;j"-R-
RRRRRRRRRRRR7_Yh7 q_hRR:1Qa)h:tR=VR"NCD#"-;-0Csk:7u1qsRFRa7zYR7qFwsR7Rq;V#NDC7:Rq _1pR
RRRRRRRRRR7RRz7aYq _1pRR:1Qa)h:tR=4R"j"jj;
--RRRRRRRRRRRRRiBpm_zaw7a_Q:)RR0LHRR:=';4'RR--BmpizVaRHRMC0HkMM8oRHOsC0MHF34R''-:RR';RjR':+RR
RRRRRRRRRRRRBmpiz_auw7a_Q:)RR0LHRR:=';4'RR--':4'R;-RR''j:
R+RRRRRRRRRRRRRiBpm_za7_pY1ua RH:RMo0CC:sR=;RjRR--j,,4.
,cRRRRRRRRRRRRRiBpmuza_Y7p_ 1auRR:HCM0oRCs:j=R;-R-R4j,,
.
RRRRRRRRRRRRRiBpm7zad)_1BRR:1Qa)h:tR=BR"pzima-";-D#CCRO08dHPR0Fkb,k0RiBpmuzaRRFsBmpizRa
RRRRRRRRRRRRBwpiA _1pRR:1Qa)h:tR=BR"pzima
";RRRRRRRRRRRRRiBpm_zaAqYu1:1RR)1aQRht:"=RV#NDC
";RRRRRRRRRRRRRiBpmuza_uAYqR11:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRpRBiamz7Y_Au1q1R1:Rah)Qt=R:RN"VD"#C;R
RRRRRRRRRRBRRpzima17_):BRR)1aQRht:"=RBmpiz;a"-C-#D0CORP8HR0Fkb,k0RpRBiamzusRFRiBpm
zaRRRRRRRRRRRRRh7Y_Q17e _1pRR:HCM0oRCs:.=RRR--..~4UM,FDC$RPRCMM
klSRRRR2RR;R
RRmRu)
a5RRRRRRRRRRRRRiBpQ:hRRRQh#_08DHFoOC_POs0F586RF0IMF2Rj;R
RRRRRRRRRRBRRpAiwRQ:Rh0R#8F_Do:HO=''j;R
RRRRRRRRRRQRRhp1 RQ:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;RRRRRRRRRRRRR1Q7 :pRRRQM#_08DHFoOC_POs0F586RF0IMF2Rj;R
RRRRRRRRRRwRRA 71pRR:Q#MR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
RRRRRRRRRRRR R)1R a:MRHR8#0_oDFH=O:';j'
RRRRRRRRRRRR R)1_ auRR:H#MR0D8_FOoH:j=''R;
RRRRRRRRRRRR)  1aR_Q:RHM#_08DHFoO':=j
';RRRRRRRRRRRRR1)  1a_RH:RM0R#8F_DoRHO:j=''R;
RRRRRRRRRRRRuq17,pw7YRR:Q#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRRRRRzR7aqY7RQ:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRRRRRRBpmiRR:mRza#_08DHFoOR;
RRRRRRRRRRRRBmpiz:aRRamzR8#0_oDFH
O;RRRRRRRRRRRRRiBpm7zaRF:Rk#0R0D8_FOoH;R
RRRRRRRRRRBRRpzima:uRR0FkR8#0_oDFH
O;RRRRRRRRRRRRRiBpm7zadRR:FRk0#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVuRpp:FRBlMbFCRM0H0#Rs;kC
-
------------------------------p-Bie7Q-------------------------B-
mmvuha hRiBp7
QeRRRRt  h)5QB
RSRR7RRQve_mR7 :aR1)tQhRR:=";."RR--",."R3"d6R",",c"R""6
RSRRtRR1h) R1:Rah)Qt=R:RN"VD"#CRR--"DVN#,C"Rs"0k
C"SRRRR
2;RRRRuam)5R
RRRRRR]RRBQpihRR:Q#hR0D8_FOoH;R
SRRRR)  1a:hRRRQh#_08DHFoOS;
RRRRRp1 d:6RRRQM#_08DHFoOS;
RRRRRiBpmRza:zRma0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRBie7QRB:RFFlbM0CMRRH#0Csk;C

MO8RFFlbM0CM#R;RR
R





