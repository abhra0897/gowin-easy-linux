`ifndef ATCIIC100_CONFIG_VH
`define ATCIIC100_CONFIG_VH
`include "ae250_config.vh"
`include "ae250_const.vh"
//	`define ATCIIC100_FIFO_DEPTH_2
//	`define ATCIIC100_FIFO_DEPTH_4
//	`define ATCIIC100_FIFO_DEPTH_8
//	`define ATCIIC100_FIFO_DEPTH_16
`endif
