--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb..4N/OGlbNbC/s#GHHDMDG/HoL/C#M_b0NsN/MdsMNl_3sIPyE84
Rf-
-
---
--
-Rl1HbRDC)RqvIEH0RM#HoRDCq)77 R11VRFsLEF0RNsC8MRN8sRIH
0C-a-RNCso0RR:XHHDM
G
DsHLNRs$HCCC;k

#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)v)h_W#RH
RRRRMoCCOsHRR5
RRRRRVRRNDlH$RR:#H0sM:oR=MR"F"MC;R
RRRRRRHRI8R0E:MRH0CCos=R:R;4jRR
RRRRRR8RN8HsI8R0E:MRH0CCos=R:R;4dRRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ERRRRRRRR80CbERR:HCM0oRCs:U=R4;g.
RRRRRRRRk8F0C_soRR:LDFFCRNM:V=RNCD#;RRRR-R-R#ENR0FkbRk0s
CoRRRRRRRR8_HMsRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#8NN0RbHMks0RCSo
RRRRs_#08NN0R#:R0MsHoS;
S_IslCF8R#:R0MsHo=R:R)"WQ_a w1Q)a
";RRRRRRRRNs88_osCRL:RFCFDN:MR=sR0kRCRRRRR-E-RNN8R8C8s#s#RCRo
RRRRR2RR;R
RRFRbs50R
RRRRRRRRz7maF:Rk#0R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRR7RRQRhR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRR7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;
RRRRRWRR :RRRRHM#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
RRRRRRRRiBpRH:RM0R#8F_Do;HORRRRR-RR-DROFRO	VRFss,NlR8N8s8,RHSM
SpmBiRR:H#MR0D8_FOoH;S
S)R1a:MRHR8#0_oDFHRO;RRRRR-R-R#sCCF0RMkRF00bkRosC
 SShRR:H#MR0D8_FOoHSRSR-C-RMHRbMVRFRFLDOs	RNSl
S
2;CRM8CHM00)$Rq_vh)
W;
ONsECH0Os0kCDRLF_O	sRNlF)VRq_vh)HWR#k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;-
-Ns00H0LkCCRoMNCs0_FssFCbsF0RVDRLF_O	sRNl:sRNO0EHCkO0sHCR#kRVMHO_M5H080Fk_osC2V;
k0MOHRFM#H0sM#o.DNP5R#:R0MsHos2RCs0kM0R#8F_Do_HOP0COFHsR#N
PsLHND#CRD:PRR8#0_oDFHPO_CFO0s'5NEEHo-DN'F8IRF0IMF2Rj;N
PsLHNDHCRRH:RMo0CC
s;LHCoMR
RVRFsHMRHR0jRFDR#PH'EoDERF
FbRRRRH5VRN'5NEEHo-RH2=4R''02RE
CMS#RRDHP52=R:R''4;C
SD
#CS#RRDHP52=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsM#;DP
8CMRs#0H.Mo#;DP
MVkOF0HMDR#P0.#soHM5:NRR8#0_oDFHPO_CFO0ss2RCs0kM0R#soHMR
H#PHNsNCLDR:#RRs#0H5MoNH'EoNE-'IDF+84RF0IMF2R4;N
PsLHNDHCRRH:RMo0CC
s;LHCoMR
RVRFsHMRHRDN'F0IRF'RNEEHoRFDFbR
RRVRHR55NH=2RR''42ER0CSM
R5R#H'-ND+FI4:2R=4R''S;
CCD#
RSR#-5HNF'DI2+4RR:=';j'
MSC8VRH;R
RCRM8DbFF;R
RskC0s#MR;M
C8DR#P0.#soHM;0
N0LsHkR0CGbO_s#FbR#:R0MsHo-;
-MOF#M0N0sR#PRND:0R#8F_Do_HOP0COFIs5HE80-84RF0IMF2RjRR:=#H0sM#o.DsP5#80_N20N;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#VOkM0MHFR0oC_FOEH_OCI0H8EH5I8R0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;N
PsLHND8CRH.Pd,HR8P,4nRP8HU8,RH,PcRP8H.8,RHRP4:MRH0CCosL;
CMoH
8RRH.PdRR:=58IH04E-2n/d;R
R84HPn=R:RH5I8-0E442/UR;
RP8HU=R:RH5I8-0E4g2/;R
R8cHPRR:=58IH04E-2;/c
8RRHRP.:5=RI0H8E2-4/
.;RHR8P:4R=IR5HE80-;42
HRRV8R5HRP4>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>.RRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8HcRR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8UHPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HnP4Rj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
R--RRHV5P8Hd>.RRRj20MEC
R--RPRRN:DR=NRPDRR+4-;
-CRRMH8RVR;
RRHV5DPNR.>R2ER0CRM
RsRRCs0kM.R5RR**PRND+RR.*5*RPRND-2Rd2R;
R#CDCR
RRCRs0MksRR5.*P*RN;D2
CRRMH8RVR;RRRRRRM
C8CRo0E_OFCHO_8IH0
E;VOkM0MHFR0oC_FOEH_OC80CbEC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLC_R8OHEFO8C_CEb0RH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0>ERRgU4.02RE
CMRRRR8E_OFCHO_b8C0:ER=nR4d;Uc
CRRDV#HRC58bR0E<U=R4Rg.NRM880CbERR>cnjgR02RE
CMRRRR8E_OFCHO_b8C0:ER=4RUg
.;RDRC#RHV5b8C0<ER=jRcgNnRM88RCEb0R.>Rj2cURC0EMR
RR_R8OHEFO8C_CEb0RR:=cnjg;R
RCHD#V8R5CEb0RR<=.UjcR8NMRb8C0>ERR.4jcRR20MEC
RRRRO8_EOFHCC_8bR0E:.=Rj;cU
CRRDV#HRC58bR0E<4=RjR.cNRM880CbERR>624.RC0EMR
RR_R8OHEFO8C_CEb0RR:=4cj.;R
RCHD#V8R5CEb0RR<=624.RC0EMR
RR_R8OHEFO8C_CEb0RR:=6;4.
CRRMH8RVR;
R0sCkRsM8E_OFCHO_b8C0
E;CRM8o_C0OHEFO8C_CEb0;k
VMHO0FoMRCI0_HE80_8lF_OU5EOFHC8_IRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDICRHE80_8lF_:URR0HMCsoC;C
Lo
HMRVRHRE5OFCHO_RI8>2RURC0EMR
RRHRI8_0El_F8U=R:RFOEH_OCI-8RRE5OFCHO_RI8lRF8U
2;RDRC#RC
RIRRHE80_8lF_:UR=EROFCHO_;I8
CRRMH8RVR;
R0sCkRsMI0H8EF_l8;_U
8CMR0oC_8IH0lE_FU8_;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=o_C0OHEFOIC_HE8058IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=nR4d/Uco_C0I0H8EF_l85_UIE_OFCHO_8IH0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CRo0E_OFCHO_b8C08E5CEb02O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=5d4nU8c/_FOEH_OC80CbE+2RR455ncdU/O8_EOFHCC_8b20ERU/R2
;
VOkM0MHFR0oC_lMk_DOCDI#58RR:HCM0o;CsOHEFOIC_8RR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCM_klODCD#RR:HCM0o;Cs
oLCHRM
RlMk_DOCD:#R=IR582-4/FOEH_OCI+8RR
4;RCRs0MksRlMk_DOCD
#;CRM8o_C0M_klODCD#
;
VOkM0MHFR0oC_x#HCM5IORR:HCM0o;CsRO8MRH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRsRRCs0kMMRIORR*8;MO
8CMR0oC_x#HC
;
VOkM0MHFR0oC_FLFD885_x#HCRR:HCM0o;CsR#I_HRxC:MRH0CCos8;R_ROI:MRH0CCosI;R_ROI:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHHM
V8R5_x#HC=R<R#I_H2xCRC0EMR
RskC0s8MR_;OI
#CDCR
RskC0sIMR_;OI
8CMR;HV
8CMR0oC_FLFD
8;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbE
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSS8E_OFCHO_8IH0RE,IE_OFCHO_8IH0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRSRRIR5HE80-/428E_OFCHO_8IH0RE,58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:R0oC_FLFDo85C#0_H5xCo_C0M_klODCD#H5I8,0ERO8_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_R8OHEFO8C_CEb02
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSRRC58b-0E482/_FOEH_OC80CbE5,R80CbE2-4/OI_EOFHCC_8b20ER4+R;
SRO#FM00NMRsxCFRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#H-I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;O#FM00NMRP#sN#D_D:PRR8#0_oDFHPO_CFO0sE5OFCHO_8IH0IE*HE80_lMk_DOCD4#-RI8FMR0Fj:2R=CRxs&FRRs#0H.Mo#5DPs_#08NN02O;
F0M#NRM0#NsPDRR:#H0sMOo5EOFHCH_I8*0EI0H8Ek_MlC_ODRD#8MFI04FR2=R:RP#D.s#0H5Mo#NsPDD_#P
2;-H-#oDMN#FRVsFRMM#-DECNb8DRLFRO	s#Nl
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,.Rd*8IH0ME_kOl_C#DD+Rd48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k.#dRF:RkL0_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRsN8C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RR--0sFRC#oH0RCs0REC#CCDO#0RHNoMDVRFRH0s#00NC-
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
RR
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjjjj"RR&Ns8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjjjjj&"RR_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjRj"&8RN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
SRDRRFNI_8R8s<"=RjjjjjjjjjRj"&8RN_osC58dRF0IMF2Rj;C
SMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjj&"RR_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjj"jjRN&R8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjj"RR&Ns8_Cno5RI8FMR0Fj
2;S8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjj"RR&Ns8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj"jjRN&R8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjRj"&8RN_osC58gRF0IMF2Rj;C
SMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDI8_N8<sR=jR"j&"RR_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDI8_N8<sR=jR''RR&Ns8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R_N8s5Co48dRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;C
SMo8RCsMCNR0Cz;46
R
RRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
R
RR8RN_osCRR<=q)77;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n114_4R
RR4RzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0SC
RORzE:	RRRHV58RN8HsI8R0E>cR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRc<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;c2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRRRRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjz.;R
RR-R-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_ncdUX:4RRLDNCHDR#1R")peq=&"RRP#sN[D5+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cXRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*d4nURc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*d4nURc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_ncdUX:4RRv)qA_4n1S4
RRRRRRRRRRRRb0FsRblNRQ575Rj2=H>RMC_so25[,7Rq7=)R>FRDI8_N84s5dFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)aS,
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7jm52>R=R0Fk_#Lk4,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;..
RRRRRRRR8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRd<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;d2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRScz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qvU.4gX:.RRLDNCHDR#1R")peq=&"RRP#sN.D5*.[+RI8FMR0F.+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gX:.RRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5UH*42g.R"&RW&"RR0HMCsoC'NHlo[C5*R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42U.4g,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*.;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gU4.RX.:qR)vnA4_
1.RRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77RR=>D_FINs885R4.8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1a
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R42=F>RkL0_k5#.H*,.[2+4,mR75Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR.<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;.2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qvcnjgX:cRRLDNCHDR#1R")peq=&"RRP#sNcD5*c[+RI8FMR0Fc+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvcnjgX:cRRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5cH*j2gnR"&RW&"RR0HMCsoC'NHlo[C5*Rc2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42cnjg,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*c;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gcjnRXc:qR)vnA4_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7R7)=D>RFNI_858s484RF0IMF2Rj,hR RR=> Rh,1R1)=)>R1Ra,
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75Rd2=F>RkL0_k5#cHc,R*d[+27,Rm25.RR=>F_k0Lck#5cH,*.[+2
,RSSSS74m52>R=R0Fk_#Lkc,5Hc+*[4R2,7jm52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>4R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF4R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR4
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq.v_jXcUURR:DCNLD#RHR)"1e=qp"RR&#NsPD*5g[R+g8MFI0gFR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUURR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*.cRU2&WR""RR&HCM0o'CsHolNC*5[g&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4.2*j,cURb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;g2
SSSLHCoMR
RRRRRRRRRRARS)_qv.UjcX:URRv)qA_4n1Sg
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7=)R>FRDI8_N84s5jFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25(RR=>F_k0LUk#5UH,*([+27,Rm25nRR=>F_k0LUk#5UH,*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75R62=F>RkL0_k5#UH*,U[2+6,mR75Rc2=F>RkL0_k5#UH*,U[2+c,mR75Rd2=F>RkL0_k5#UH*,U[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.=2R>kRF0k_L#HU5,[U*+,.2R57m4=2R>kRF0k_L#HU5,[U*+,42R57mj=2R>kRF0k_L#HU5,[U*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRQR7u25jRR=>HsM_Cgo5*U[+27,Rmju52>R=RsbNH_0$LUk#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>42jRRMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R24jRR<=Ns8_CNo58I8sHE80-84RF0IMFjR42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcSzjRR:H5VRNs88I0H8ERR>4Rj2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_4.4cXnRR:DCNLD#RHR)"1e=qp"RR&#NsPDU54*4[+UFR8IFM0R*4U[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXnRR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*4.Rc2&WR""RR&HCM0o'CsHolNC*5[4RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424cj.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+2U*42S;
SCSLo
HMRRRRRRRRRRRRSqA)vj_4.4cXnRR:)Aqv41n_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7=)R>FRDI8_N8gs5RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,RR
RRRRRRRRRRRRRRRRRRRRRRRRRWRR >R=R0Is_5CMHR2,BRpi=B>RpRi,74m56=2R>kRF0k_L#54nHn,4*4[+6R2,74m5c=2R>kRF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4Rd2=F>RkL0_kn#454H,n+*[4,d2R57m4R.2=F>RkL0_kn#454H,n+*[4,.2R57m4R42=F>RkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7524jRR=>F_k0L4k#n,5H4[n*+24j,mR75Rg2=F>RkL0_kn#454H,n+*[gR2,7Um52>R=R0Fk_#Lk4Hn5,*4n[2+U,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR75R(2=F>RkL0_kn#454H,n+*[(R2,7nm52>R=R0Fk_#Lk4Hn5,*4n[2+n,mR75R62=F>RkL0_kn#454H,n+*[6
2,SRSSR7RRm25cRR=>F_k0L4k#n,5H4[n*+,c2R57md=2R>kRF0k_L#54nHn,4*d[+27,Rm25.RR=>F_k0L4k#n,5H4[n*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4=2R>kRF0k_L#54nHn,4*4[+27,Rm25jRR=>F_k0L4k#n,5H4[n*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_soU54*4[+(FR8IFM0R*4U[n+42R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4u52>R=RsbNH_0$L4k#n,5H.+*[4R2,75muj=2R>NRbs$H0_#Lk4Hn5,[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co4[U*2=R<R0Fk_#Lk4Hn5,*4n[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R42<F=RkL0_kn#454H,n+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R.2<F=RkL0_kn#454H,n+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rd2<F=RkL0_kn#454H,n+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rc2<F=RkL0_kn#454H,n+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R62<F=RkL0_kn#454H,n+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rn2<F=RkL0_kn#454H,n+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R(2<F=RkL0_kn#454H,n+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+RU2<F=RkL0_kn#454H,n+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rg2<F=RkL0_kn#454H,n+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24jRR<=F_k0L4k#n,5H4[n*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+4<2R=kRF0k_L#54nHn,4*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24.RR<=F_k0L4k#n,5H4[n*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+d<2R=kRF0k_L#54nHn,4*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24cRR<=F_k0L4k#n,5H4[n*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+6<2R=kRF0k_L#54nHn,4*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24nRR<=bHNs0L$_kn#45.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[(+42=R<RsbNH_0$L4k#n,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d
cSzdRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>gRR2oCCMsCN0
RSRRORzDR	:bOsFCR##5iBp2S
SRCRLo
HMSRSRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRRRRNRR8osC58N8s8IH04E-RI8FMR0Fg<2R=8RN_osC58N8s8IH04E-RI8FMR0Fg
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	S;
RRRRzRcc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzRc6:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SS8CMRMoCC0sNCcRz6S;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSSc:nRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0Rnzc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSSc:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qv6X4.d:.RRLDNCHDR#1R")peq=&"RRP#sNdD5n+*[d8nRF0IMFnRd*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.RR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCH4*6.&2RR""WRH&RMo0CCHs'lCNo5d[*n&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+462*4R.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42d;n2
SSSLHCoMR
RRRRRRRRRRRRRRRRRRRRRRRRRAv)q_.64XRd.:qR)vnA4_n1d
RRRRRRRRRRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Cod[n*+Rd48MFI0dFRn2*[,7Rq7=)R>IDF_8N8sR5U8MFI0jFR2 ,Rh>R=R, hR)11RR=>),1a
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRWRR >R=R0Is_5CMHR2,BRpi=B>RpRi,7dm54=2R>kRF0k_L#5d.H.,d*d[+4R2,7dm5j=2R>kRF0k_L#5d.H.,d*d[+j
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.gRR=>F_k0Ldk#.,5Hd[.*+2.g,mR752.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR752.(RR=>F_k0Ldk#.,5Hd[.*+2.(,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5n=2R>kRF0k_L#5d.H.,d*.[+nR2,7.m56=2R>kRF0k_L#5d.H.,d*.[+6R2,7.m5c=2R>kRF0k_L#5d.H.,d*.[+c
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR752..RR=>F_k0Ldk#.,5Hd[.*+2..,mR752.4RR=>F_k0Ldk#.,5Hd[.*+2.4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5j=2R>kRF0k_L#5d.H.,d*.[+jR2,74m5g=2R>kRF0k_L#5d.H.,d*4[+gR2,74m5U=2R>kRF0k_L#5d.H.,d*4[+U
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7524(RR=>F_k0Ldk#.,5Hd[.*+24(,mR7524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR75246RR=>F_k0Ldk#.,5Hd[.*+246,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR74m5c=2R>kRF0k_L#5d.H.,d*4[+cR2,74m5d=2R>kRF0k_L#5d.H.,d*4[+dR2,74m5.=2R>kRF0k_L#5d.H.,d*4[+.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4542>R=R0Fk_#LkdH.5,*d.[4+427,Rmj542>R=R0Fk_#LkdH.5,*d.[j+427,Rm25gRR=>F_k0Ldk#.,5Hd[.*+,g2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Um52>R=R0Fk_#LkdH.5,*d.[2+U,mR75R(2=F>RkL0_k.#d5dH,.+*[(R2,7nm52>R=R0Fk_#LkdH.5,*d.[2+n,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m6=2R>kRF0k_L#5d.H.,d*6[+27,Rm25cRR=>F_k0Ldk#.,5Hd[.*+,c2R57md=2R>kRF0k_L#5d.H.,d*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75R.2=F>RkL0_k.#d5dH,.+*[.R2,74m52>R=R0Fk_#LkdH.5,*d.[2+4,mR75Rj2=F>RkL0_k.#d5dH,.2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u25dRR=>bHNs0L$_k.#d5cH,*d[+27,Rm.u52>R=RsbNH_0$Ldk#.,5Hc+*[.
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_k.#d5cH,*4[+27,Rmju52>R=RsbNH_0$Ldk#.,5Hc2*[2R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4<2R=kRF0k_L#5d.H.,d*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[d<2R=kRF0k_L#5d.H.,d*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[6<2R=kRF0k_L#5d.H.,d*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[(<2R=kRF0k_L#5d.H.,d*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[g<2R=kRF0k_L#5d.H.,d*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+42=R<R0Fk_#LkdH.5,*d.[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+42=R<R0Fk_#LkdH.5,*d.[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+42=R<R0Fk_#LkdH.5,*d.[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+42=R<R0Fk_#LkdH.5,*d.[(+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+42=R<R0Fk_#LkdH.5,*d.[g+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+.2=R<R0Fk_#LkdH.5,*d.[4+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[d+.2=R<R0Fk_#LkdH.5,*d.[d+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+.2=R<R0Fk_#LkdH.5,*d.[6+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[(+.2=R<R0Fk_#LkdH.5,*d.[(+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[g+.2=R<R0Fk_#LkdH.5,*d.[g+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[4+d2=R<R0Fk_#LkdH.5,*d.[4+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2ddRR<=bHNs0L$_k.#d5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+6<2R=NRbs$H0_#LkdH.5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSCRM8oCCMsCN0R(zc;S
SCRM8oCCMsCN0Rczc;C
SMo8RCsMCNR0Cz;cd
M
C8sRNO0EHCkO0sLCRD	FO_lsN;N

sHOE00COkRsCMsF_IE_OCRO	F)VRq_vh)HWR#k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kMh5"FCRsNI8/sCH0RMOFVODH0EROC3O	Rl1Hk0DNHRFMllH#NE0OR#bF#DHLC!R!"
2;RDRC#RC
RsRRCs0kM'5"MsF_IE_OC'O	RRH#0REC#CNlRRN#'FLDOs	_NRl'VRFs#oHMDbCRFRs0)#qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
0N0skHL0oCRCsMCNs0F_bsCFRs0:0R#soHM;-
-Ns00H0LkCCRoMNCs0_FssFCbsF0RVFRM__sIOOEC	RR:NEsOHO0C0CksRRH#VOkM_HHM085N8ss_C;o2
MVkOF0HM0R#soHM.P#D5:NRRs#0H2MoR0sCkRsM#_08DHFoOC_POs0FR
H#PHNsNCLDRP#DR#:R0D8_FOoH_OPC05FsNH'EoNE-'IDFRI8FMR0Fj
2;PHNsNCLDR:HRR0HMCsoC;C
Lo
HMRFRVsRRHHjMRRR0F#'DPEEHoRFDFbR
RRVRHR55NNH'EoHE-2RR='24'RC0EMR
SRP#D5RH2:'=R4
';S#CDCR
SRP#D5RH2:'=Rj
';S8CMR;HV
CRRMD8RF;Fb
sRRCs0kMDR#PC;
M#8R0MsHoD.#PV;
k0MOHRFM#.DP#H0sMNo5R#:R0D8_FOoH_OPC02FsR0sCkRsM#H0sMHoR#N
PsLHND#CRR#:R0MsHo'5NEEHo-DN'F4I+RI8FMR0F4
2;PHNsNCLDR:HRR0HMCsoC;C
Lo
HMRFRVsRRHHNMR'IDFRR0FNH'EoDERF
FbRRRRH5VRN25HR'=R4R'20MEC
RSR#-5HNF'DI2+4RR:=';4'
DSC#SC
R5R#H'-ND+FI4:2R=jR''S;
CRM8H
V;RMRC8FRDF
b;RCRs0MksR
#;CRM8#.DP#H0sM
o;Ns00H0LkCORG_Fbsb:#RRs#0H;Mo
O--F0M#NRM0#NsPDRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0Fj:2R=0R#soHM.P#D50s#_08NN
2;-L-RCMoHRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#k
VMHO0FoMRCO0_EOFHCH_I850EI0H8ERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;PHNsNCLDRP8HdR.,84HPn8,RH,PURP8Hc8,RH,P.RP8H4RR:HCM0o;Cs
oLCHRM
RP8Hd:.R=IR5HE80-/42d
n;RHR8PR4n:5=RI0H8E2-4/;4U
8RRHRPU:5=RI0H8E2-4/
g;RHR8P:cR=IR5HE80-/42cR;
RP8H.=R:RH5I8-0E4.2/;R
R84HPRR:=58IH04E-2R;
RRHV5P8H4RR>j02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RH5VR8.HPRj>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
HRRV8R5HRPc>2RjRC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RVRHRH58P>URRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
RRHV5P8H4>nRRRj20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RV-;
-HRRV8R5H.PdRj>R2ER0C-M
-RRRRDPNRR:=PRND+;R4
R--R8CMR;HV
HRRVPR5N>DRRR.20MECRR
RRCRs0MksRR5.*P*RN+DRR*.R*PR5N-DRR2d2;R
RCCD#
RRRR0sCkRsM5*.R*NRPD
2;RMRC8VRH;M
C8CRo0E_OFCHO_8IH0
E;VOkM0MHFR0oC_FOEH_OC80CbEC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLC_R8OHEFO8C_CEb0RH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0>ERRgU4.02RE
CMRRRR8E_OFCHO_b8C0:ER=nR4d;Uc
CRRDV#HRC58bR0E<U=R4Rg.NRM880CbERR>cnjgR02RE
CMRRRR8E_OFCHO_b8C0:ER=4RUg
.;RDRC#RHV5b8C0<ER=jRcgNnRM88RCEb0R.>Rj2cURC0EMR
RR_R8OHEFO8C_CEb0RR:=cnjg;R
RCHD#V8R5CEb0RR<=.UjcR8NMRb8C0>ERR.4jcRR20MEC
RRRRO8_EOFHCC_8bR0E:.=Rj;cU
CRRDV#HRC58bR0E<4=RjR.cNRM880CbERR>624.RC0EMR
RR_R8OHEFO8C_CEb0RR:=4cj.;R
RCHD#V8R5CEb0RR<=624.RC0EMR
RR_R8OHEFO8C_CEb0RR:=6;4.
CRRMH8RVR;
R0sCkRsM8E_OFCHO_b8C0
E;CRM8o_C0OHEFO8C_CEb0;k
VMHO0FoMRCI0_HE80_8lF_OU5EOFHC8_IRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDICRHE80_8lF_:URR0HMCsoC;C
Lo
HMRVRHRE5OFCHO_RI8>2RURC0EMR
RRHRI8_0El_F8U=R:RFOEH_OCI-8RRE5OFCHO_RI8lRF8U
2;RDRC#RC
RIRRHE80_8lF_:UR=EROFCHO_;I8
CRRMH8RVR;
R0sCkRsMI0H8EF_l8;_U
8CMR0oC_8IH0lE_FU8_;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=o_C0OHEFOIC_HE8058IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=nR4d/Uco_C0I0H8EF_l85_UIE_OFCHO_8IH0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CRo0E_OFCHO_b8C08E5CEb02O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=5d4nU8c/_FOEH_OC80CbE+2RR455ncdU/O8_EOFHCC_8b20ERU/R2
;
VOkM0MHFR0oC_lMk_DOCDI#58RR:HCM0o;CsOHEFOIC_8RR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCM_klODCD#RR:HCM0o;Cs
oLCHRM
RlMk_DOCD:#R=IR582-4/FOEH_OCI+8RR
4;RCRs0MksRlMk_DOCD
#;CRM8o_C0M_klODCD#
;
VOkM0MHFR0oC_x#HCM5IORR:HCM0o;CsRO8MRH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRsRRCs0kMMRIORR*8;MO
8CMR0oC_x#HC
;
VOkM0MHFR0oC_FLFD885_x#HCRR:HCM0o;CsR#I_HRxC:MRH0CCos8;R_ROI:MRH0CCosI;R_ROI:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHHM
V8R5_x#HC=R<R#I_H2xCRC0EMR
RskC0s8MR_;OI
#CDCR
RskC0sIMR_;OI
8CMR;HV
8CMR0oC_FLFD
8;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbE
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSS8E_OFCHO_8IH0RE,IE_OFCHO_8IH0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:o=RCL0_F8FD50oC_x#HCC5o0k_MlC_OD5D#I0H8E8,R_FOEH_OCI0H8Eo2,CM0_kOl_C#DD5b8C0RE,8E_OFCHO_b8C02E2,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRo0H_#xoC5CM0_kOl_C#DD58IH0RE,IE_OFCHO_8IH0,E2o_C0M_klODCD#C58b,0EROI_EOFHCC_8b20E2S,
SSSSSSSSSRSRRIR5HE80-/428E_OFCHO_8IH0RE,58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:R0oC_FLFDo85C#0_H5xCo_C0M_klODCD#H5I8,0ERO8_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_R8OHEFO8C_CEb02
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRRC#0_H5xCo_C0M_klODCD#H5I8,0EROI_EOFHCH_I820E,0oC_lMk_DOCD8#5CEb0,_RIOHEFO8C_CEb02
2,SSSSSSSSSRSRRC58b-0E482/_FOEH_OC80CbE5,R80CbE2-4/OI_EOFHCC_8b20ER4+R;
SRO#FM00NMRsxCFRR:#_08DHFoOC_POs0F5FOEH_OCI0H8EH*I8_0EM_klODCD#H-I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;O#FM00NMRP#sN#D_D:PRR8#0_oDFHPO_CFO0sE5OFCHO_8IH0IE*HE80_lMk_DOCD4#-RI8FMR0Fj:2R=CRxs&FRRs#0H.Mo#5DPs_#08NN02O;
F0M#NRM0#NsPDRR:#H0sMOo5EOFHCH_I8*0EI0H8Ek_MlC_ODRD#8MFI04FR2=R:RP#D.s#0H5Mo#NsPDD_#P
2;-H-#oDMN#FRVsFRMM#-DECNb8DRLFRO	s#Nl
b0$CkRF0k_L#04_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#4:kRF0k_L#04_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0c_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkcRR:F_k0Lck#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kR#U:NRbs$H0_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,dI.*HE80_lMk_DOCDd#+4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lkd:.RR0Fk_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRsN8C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RR--0sFRC#oH0RCs0REC#CCDO#0RHNoMDVRFRH0s#00NC-
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
RR
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjjjj"RR&Ns8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjjjjj&"RR_N8s5Co4FR8IFM0R;j2
MSC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRRd2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjjRj"&8RN_osC58.RF0IMF2Rj;C
SMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
SRDRRFNI_8R8s<"=RjjjjjjjjjRj"&8RN_osC58dRF0IMF2Rj;C
SMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjj&"RR_N8s5CocFR8IFM0R;j2
MSC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjj"jjRN&R8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjj"RR&Ns8_Cno5RI8FMR0Fj
2;S8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjj"RR&Ns8_C(o5RI8FMR0Fj
2;S8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj"jjRN&R8C_soR5U8MFI0jFR2S;
CRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjRj"&8RN_osC58gRF0IMF2Rj;C
SMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co48jRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RSRRFRDI8_N8<sR=jR"j&"RR_N8s5Co484RF0IMF2Rj;C
SMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RSRRFRDI8_N8<sR=jR''RR&Ns8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R_N8s5Co48dRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;C
SMo8RCsMCNR0Cz;46
R
RRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
R
RR8RN_osCRR<=q)77;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n114_4R
RR4RzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0SC
RORzE:	RRRHV58RN8HsI8R0E>cR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRc<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;c2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRRRRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjz.;R
RR-R-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRR.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_ncdUX:4RRLDNCHDR#1R")peq=&"RRP#sN[D5+R42&,R"RQW)av _m=7 "RR&Ils_F;8C
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cXRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*d4nURc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*d4nURc,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_ncdUX:4RRv)qA_4n1S4
RRRRRRRRRRRRb0FsRblNRQ575Rj2=H>RMC_so25[,7Rq7=)R>FRDI8_N84s5dFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)aS,
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7jm52>R=R0Fk_#Lk4,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;..
RRRRRRRR8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRd<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;d2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRScz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rd2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.6:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCS
SS0N0skHL0GCROs_bFRb#FAVR)_qvU.4gX:.RRLDNCHDR#1R")peq=&"RRP#sN.D5*.[+RI8FMR0F.+*[4&2RRR",Wa)Q m_v7" =RI&RsF_l8
C;RRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gX:.RRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5UH*42g.R"&RW&"RR0HMCsoC'NHlo[C5*R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*42U.4g,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*.;S
SSoLCHRM
RRRRRRRRRSRRAv)q_gU4.RX.:qR)vnA4_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7R7)=D>RFNI_858s48.RF0IMF2Rj,hR RR=> Rh,1R1)=)>R1
a,SSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4=2R>kRF0k_L#H.5,[.*+,42R57mj=2R>kRF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5[.*2=R<R0Fk_#Lk.,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5.[2+4RR<=F_k0L.k#5.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(z.;R
RRSRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RS

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHR85N8HsI8R0E>.R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF.R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR.
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAqcv_jXgncRR:DCNLD#RHR)"1e=qp"RR&#NsPD*5c[R+c8MFI0cFR*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqcv_jXgncRR:DCNLD#RHR1"Aa&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHj*cgRn2&WR""RR&HCM0o'CsHolNC*5[c&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5HRR+4c2*j,gnRb8C02E2R"&RX&"RR0HMCsoC'NHlo5C5[2+4*;c2
SSSLHCoMR
RRRRRRRRRRARS)_qvcnjgX:cRRv)qA_4n1Sc
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7=)R>FRDI8_N84s54FR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57md=2R>kRF0k_L#Hc5,*Rc[2+d,mR75R.2=F>RkL0_k5#cH*,c[2+.,SR
S7SSm254RR=>F_k0Lck#5cH,*4[+27,Rm25jRR=>F_k0Lck#5RH,c2*[2R;
RRRRRRRRRRRRRFRRks0_Cco5*R[2<F=RkL0_k5#cH*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[4<2R=kRF0k_L#Hc5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R.2<F=RkL0_k5#cH*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+dRR<=F_k0Lck#5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.zd;R
RRSRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR244RMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R244RR<=Ns8_CNo58I8sHE80-84RF0IMF4R42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRSd:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSNSS0H0sLCk0R_GObbsF#VRFRqA)vj_.cUUXRD:RNDLCRRH#"e1)q"p=R#&RsDPN5[g*+8gRF0IMF*Rg[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUXRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*c.jU&2RR""WRH&RMo0CCHs'lCNo5g[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2j*.cRU,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42g
2;SLSSCMoH
RRRRRRRRRRRR)SAq.v_jXcUURR:)Aqv41n_gR
SRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)>R=RIDF_8N8sj54RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7(m52>R=R0Fk_#LkU,5HU+*[(R2,7nm52>R=R0Fk_#LkU,5HU+*[nR2,
SSSS57m6=2R>kRF0k_L#HU5,[U*+,62R57mc=2R>kRF0k_L#HU5,[U*+,c2R57md=2R>kRF0k_L#HU5,[U*+,d2RS
SSmS75R.2=F>RkL0_k5#UH*,U[2+.,mR75R42=F>RkL0_k5#UH*,U[2+4,mR75Rj2=F>RkL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQju52>R=R_HMs5Cog+*[UR2,75muj=2R>NRbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
(;RRRRRMSC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1Uz
Sd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERRR4j2CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFjR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRj
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RjM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq4v_jX.c4:nRRLDNCHDR#1R")peq=&"RRP#sN4D5U+*[48URF0IMFUR4*4[+2RR&"W,R) Qa_7vm R="&sRI_8lFCR;
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4:nRRLDNCHDR#AR"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*j2.cR"&RW&"RR0HMCsoC'NHlo[C5*24UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05R5H+2R4*.4jc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[442*U
2;SLSSCMoH
RRRRRRRRRRRR)SAq4v_jX.c4:nRRv)qA_4n1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7R7)=D>RFNI_858sgFR8IFM0R,j2RR h= >Rh1,R1=)R>1R)a
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4R62=F>RkL0_kn#454H,n+*[4,62R57m4Rc2=F>RkL0_kn#454H,n+*[4,c2RS
SSmS7524dRR=>F_k0L4k#n,5H4[n*+24d,mR7524.RR=>F_k0L4k#n,5H4[n*+24.,mR75244RR=>F_k0L4k#n,5H4[n*+244,SR
S7SSmj542>R=R0Fk_#Lk4Hn5,*4n[j+427,Rm25gRR=>F_k0L4k#n,5H4[n*+,g2R57mU=2R>kRF0k_L#54nHn,4*U[+2S,
S7SSm25(RR=>F_k0L4k#n,5H4[n*+,(2R57mn=2R>kRF0k_L#54nHn,4*n[+27,Rm256RR=>F_k0L4k#n,5H4[n*+,62
SSSRRRR7cm52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR75Rd2=F>RkL0_kn#454H,n+*[dR2,7.m52>R=R0Fk_#Lk4Hn5,*4n[2+.,S
SRRRRRRRR74m52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR75Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ=uR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_kn#45.H,*4[+27,Rmju52>R=RsbNH_0$L4k#n,5H.2*[2R;
RRRRRRRRRRRRRFRRks0_C4o5U2*[RR<=F_k0L4k#n,5H4[n*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4<2R=kRF0k_L#54nHn,4*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[.<2R=kRF0k_L#54nHn,4*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[d<2R=kRF0k_L#54nHn,4*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[c<2R=kRF0k_L#54nHn,4*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[6<2R=kRF0k_L#54nHn,4*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[n<2R=kRF0k_L#54nHn,4*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[(<2R=kRF0k_L#54nHn,4*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[U<2R=kRF0k_L#54nHn,4*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[g<2R=kRF0k_L#54nHn,4*g[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rj2<F=RkL0_kn#454H,n+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[4+42=R<R0Fk_#Lk4Hn5,*4n[4+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R.2<F=RkL0_kn#454H,n+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[d+42=R<R0Fk_#Lk4Hn5,*4n[d+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rc2<F=RkL0_kn#454H,n+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[6+42=R<R0Fk_#Lk4Hn5,*4n[6+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rn2<b=RN0sH$k_L#54nH*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24(RR<=bHNs0L$_kn#45.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.zc;R
RRSRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1
dnSdzcRH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80Rg>RRo2RCsMCN
0CSRRRRDzO	b:RsCFO#5#RB2pi
RSSRoLCHSM
SRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMS
SRRRRR8RNs5CoNs88I0H8ER-48MFI0gFR2=R<R_N8s5CoNs88I0H8ER-48MFI0gFR2S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
SRzRRc:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>2RgRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HOSzSSc:6RRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SISSsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSCRM8oCCMsCN0R6zc;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSznRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0Cz;cn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCS#
ScSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
SSSNs00H0LkCORG_FbsbF#RV)RAq6v_4d.X.RR:DCNLD#RHR)"1e=qp"RR&#NsPDn5d*d[+nFR8IFM0R*dn[2+4R"&R,)RWQ_a v m7=&"RR_IslCF8;R
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..XdRD:RNDLCRRH#"aA1"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*.642RR&"RW"&MRH0CCosl'HN5oC[n*d2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R24*6.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4d2*n
2;SLSSCMoH
SSSSqA)v4_6..XdR):Rq4vAnd_1nR
RRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7R7)=F>DI8_N8Us5RI8FMR0FjR2, =hR>hR ,1R1)>R=Ra)1,S
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm45d2>R=R0Fk_#LkdH.5,*d.[4+d27,Rmj5d2>R=R0Fk_#LkdH.5,*d.[j+d2S,
S7SSmg5.2>R=R0Fk_#LkdH.5,*d.[g+.27,RmU5.2>R=R0Fk_#LkdH.5,*d.[U+.27,Rm(5.2>R=R0Fk_#LkdH.5,*d.[(+.2S,
S7SSmn5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rmc5.2>R=R0Fk_#LkdH.5,*d.[c+.2S,
S7SSmd5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.5.2>R=R0Fk_#LkdH.5,*d.[.+.27,Rm45.2>R=R0Fk_#LkdH.5,*d.[4+.2S,
S7SSmj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rmg542>R=R0Fk_#LkdH.5,*d.[g+427,RmU542>R=R0Fk_#LkdH.5,*d.[U+42S,
S7SSm(542>R=R0Fk_#LkdH.5,*d.[(+427,Rmn542>R=R0Fk_#LkdH.5,*d.[n+427,Rm6542>R=R0Fk_#LkdH.5,*d.[6+42S,
S7SSmc542>R=R0Fk_#LkdH.5,*d.[c+427,Rmd542>R=R0Fk_#LkdH.5,*d.[d+427,Rm.542>R=R0Fk_#LkdH.5,*d.[.+42
,RSSSS74m54=2R>kRF0k_L#5d.H.,d*4[+4R2,74m5j=2R>kRF0k_L#5d.H.,d*4[+jR2,7gm52>R=R0Fk_#LkdH.5,*d.[2+g,SR
S7SSm25URR=>F_k0Ldk#.,5Hd[.*+,U2R57m(=2R>kRF0k_L#5d.H.,d*([+27,Rm25nRR=>F_k0Ldk#.,5Hd[.*+,n2RS
SSmS75R62=F>RkL0_k.#d5dH,.+*[6R2,7cm52>R=R0Fk_#LkdH.5,*d.[2+c,mR75Rd2=F>RkL0_k.#d5dH,.+*[dR2,
SSSS57m.=2R>kRF0k_L#5d.H.,d*.[+27,Rm254RR=>F_k0Ldk#.,5Hd[.*+,42R57mj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5Rd2=b>RN0sH$k_L#5d.H*,c[2+d,mR7u25.RR=>bHNs0L$_k.#d5cH,*.[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5R42=b>RN0sH$k_L#5d.H*,c[2+4,mR7u25jRR=>bHNs0L$_k.#d5cH,*2[2;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SCSSMo8RCsMCNR0Cz;c(
CSSMo8RCsMCNR0Cz;cc
MSC8CRoMNCs0zCRc
d;
8CMRONsECH0Os0kCFRM__sIOOEC	
;
-p-RNR#0HDlbCMlC0HN0FHMR#CR8VDNk0s
NO0EHCkO0s#CRCODC0N_slVRFRv)qhW_)R
H#VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEO;
F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8RO#FM00NMRVDC0P_FC:sRR0HMCsoCRR:=5855CEb0R4+R6l2RFd8R./2RR24n;RRRRRRRRRRRRRRRRRRRRRRRR-R-RFyRVqR)vX4n4M1RCCC88FRVsCRDVF0RPRCsI8Fs#$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_ODRD#8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COFcs5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
R
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"j"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<=""jjRN&R8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR''RR&Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
RRRRRzcRH:RVNR58I8sHE80Rc>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<N=R8C_soR5c8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
c;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR6R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
6;RRRRzRnR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR(:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRRRRRCRM8oCCMsCN0R;z(
RRRRRzURH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_soR;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RRgRzRRR:H5VRNs88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRNRR8C_so=R<R7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4:jRRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4Rz4RR:VRFsHMRHRk5MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4.:VRHR85N8HsI8R0E>2R6RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5_N8s5CoNs88I0H8ER-48MFI06FR2RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RR62=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4.
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz4RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4RzcRR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*2d.R"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEH55R4+R2.*d,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRv)qd4.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CHM52W,RBRpi=B>RpRi,m>R=R0Fk_#Lk5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0Rcz4;R
RRRRRRMRC8CRoMNCs0zCR4R4;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR6z4RH:RVDR5C_V0FsPCR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR4n:VRHR85N8HsI8R0E>2R6RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDR#2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R6RM=RkOl_C#DD2MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4n
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRR(z4RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4(
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CRRRRRRRRzR4U:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCDd#*.&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC58b20ER"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=R0Fk_#Lk5lMk_DOCD[#,2
2;RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#k5MlC_OD,D#[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0RUz4;R
RRRRRRMRC8CRoMNCs0zCR4R6;RRRRRRRRRC

MN8RsHOE00COkRsC#CCDOs0_N
l;
