@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ua_)mmu1QQam;h"
R
R`OHMDCk8R0"#8P_FDN_0#E	3"`

HCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0M`C
CHM8V/R/m_epQahQ_tv1
H
`VV8CRpme_1q1 _)am
h
RDRNI#N$R5@@`pme_1)  1a_QqthpsRFR#0C0G_CbRs2LHCoMR
RRVRHRm5`e)p_ a1 _t1QhRqp!4=R'2LjRoLCHRM
RRRRRqq_1)1 a)_um1umQmaQh:_uR#N#CRs05#0C0G_Cb!sR='R4LRj2CCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHRpwq12 ";R
RRMRC8R
RCRM8/N/RD$IN#`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#C
RRRRNRRD$IN#@R@5e`mp _)1_ a1hQtqFpRs0R5C_#0CsGbR0^RC_#0CsGb2L2RCMoH
RRRRRRRRRHV5e`mp _)1_ a1hQtq!pR='R4LRj2
RRRRRRRRLRRCMoH
RRRRRRRRRRRRqq_1)1 a)_um1umQmaQhZ_X__mhaa 1_Ru:
RRRRRRRRRRRR#N#CRs0555!fkH#MF	MI0M5C_#0CsGb2R22=4=R'2L4
RRRRRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RRRRRRRRRMRC8R
RRRRRCRM8/N/RD$IN#R

RM`C8RHV/m/ReQp_vQupB_QaX B]Bmi_w
w
`8CMH/VR/eRmpB_X]i B_wmw
C
`MV8HRR//m_epq 11)ma_h



