@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)aa_)1qhQmaQh
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_qa)ha1QQ_mhuR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RC50#C0_GRbs=#=R00Ns_N#00RC2|R=>50R5C_#0CsGbRR==f#bN005#N_s0#00NCR22|R|
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0R5C_#0CsGbRR==f#bN0C5MG#0_0CN0222R;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_qa)ha1QQ_mhXmZ_h _a1 a_X_u)uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R5RR!H5f#	kMMMFI5#0C0G_Cb2s22R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aah)q1QQamXh_Zh_m_q1a)1a_a qa_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5f!5HM#k	IMFM05#N_s0#00NC222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)aa_)1qhQmaQhZ_X__mhha X_q1aau _;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RR0R5C_#0CsGbRR==#s0N00_#N20CR>|-R55!fkH#MF	MIMM5C_G0#00NC222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )_qa)ha1QQ_mhuN:R#s#C0sRbFsbC05$Rq 11)aa_)1qhQmaQh2_u
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HMsR0NHM#0MHFCV8RsRFlPkNDC0R#N_s0#00NCFR0RPNRNCDkREF0C0sRERNMM0CG_N#002C";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 a)_aqQh1ahQm__XZmah_ _1a )Xu_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a)_aqQh1ahQm__XZmah_ _1a )Xu_
u2RRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
R
RRRRRR_Rqq 11)aa_)1qhQmaQhZ_X__mh1)aqaa_1q_a uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_qa)ha1QQ_mhXmZ_ha_1q_)a1aaq 2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N#0s#0_0CN0RMOF0MNH#RRXFZsR"
2;
RRRRRRRRqq_1)1 a)_aqQh1ahQm__XZmhh_ _Xa1aaq :_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)aa_)1qhQmaQhZ_X__mhha X_q1aau _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"MG#0_0CN0RMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w

R
RRRRRC
M8RRRRRmR`eqp_1v1z RR:LHCoMRR:F_PDNk##lRC
RRRRRvRR_1q1 _)aah)q1QQamuh_:#RN#CklRFbsb0Cs$qR51)1 a)_aqQh1ahQm_;u2
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )_qa)ha1QQ_mhXmZ_h _a1 a_X_u)uR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qa)ha1QQ_mhXmZ_h _a1 a_X_u)u
2;
RRRRRRRRqv_1)1 a)_aqQh1ahQm__XZm1h_aaq)_q1aau _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aah)q1QQamXh_Zh_m_q1a)1a_a qa_;u2
R
RRRRRR_Rvq 11)aa_)1qhQmaQhZ_X__mhha X_q1aau _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aah)q1QQamXh_Zh_m_Xh aa_1q_a u
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
V`H8RCVm_epB me)h_m
C
oMNCs0
C
RRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RH5VRm_epB me)q_A1_QBmRh2LHCoMRR:F_PDOCFPsN_L#
HO
RRROCFPs0_#N_s0#00NCR:
RFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRC50#C0_GRbs=#=R00Ns_N#002C2RR2
RRRRRRRRRRRRRRRRRDFP_POFC0s_50"#N_s0#00NCFROPCCs8;"2
CRRM
8
R8CM
M
C8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



