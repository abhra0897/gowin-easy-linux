
@ER--=========m==F=FF=========================================FmFF========-
-RR=RB$FbsEHo0BR52jR.4.c-jR4(tHFIMCR1lFHOMO8k0RFsaECOMFFDoB$RFp3,0
83-=-RRRRRRRRRRRRRRRRRRRRRRDqDRosHER0#sCC#s8PC3-
-R====================================================================-=
--
-R_R_RRRRR_R_RRRRR_R_
R--R\\RRRRR/\RRRRRR/RR/RwRrHRDCMCNlR9RRRHbsl$_#ME3P8-
-R\RRRR\R/\R/RR\R/RR/RrRR7OC#s0HbHRFM9WRt.eqR]R7pVOkM0MHFN#DR$EM0C##HRLDHs$Ns
R--R\RRRR\//\RRRR\//RRRRaRrH#lC0bNlR9RRRCakRsqbH.DR6cR4::jjd.jRj
4(-R-RR\RRRRR/R\RRRRR/RRRRRCrPsF#HMRRRRRR9433(n-
-RRRRR/R\RRRRR/R\RRRRR
RR---
-=R==========FmFF========================================m==F=FF=====
==
-
--------------------------ObN	CNoRFoDL-ND-----------------------------p

QqA))HYRC;CCR1
z CRHC#C30D8_FOoH_n44cD3ND
;RkR#CQ   371a_tpmQqB_)]Qa3pqp;#
kC RQ 1 3ap7_mBtQ_1zhQ th7p3qp
;
uiqBqRt ObFlFMMC0Q#R1RR
R0RN0LsHkR0C#_$MLODN	F_LGL:RFCFDN;MR
RRRNs00H0LkC$R#MD_LN_O	LRFGFBVRFFlbM0CM#RR:b	NONRoCH0#Rs;kC
RRRNs00H0LkCDRLN_O	L_FGb_N8b:HMRs#0H;Mo
RRRNs00H0LkC$R#MF_MbMskCRR:LDFFC;NM
RRRNs00H0LkCORG_blN:0R#soHM;R
RR0N0skHL0GCRON_lbVRFRlBFbCFMMR0#:NRbOo	NC#RHRk"D0R";S-
-b	NONRoCoRDLH-#
-HS#oDMNR)t1hRR:#_08DHFoO=R:R''4;-
-CRM8o;DL
b--NNO	oLCRFR8$oRDL
C--Mo8RD
L;-----------------------------1-t)---------------------------------------
m
Bvhum RhatR1)
RRRR)uma
R5RRRRRRRRR)t1QRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVtR1):FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0#CR$MM_FkbsMFCRV1Rt)RR:BbFlFMMC0#RHRk0sC-;
-------------------------apz4----------------------------
--Bumvmhh azRpa
4RRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"Rj"2R;
RuRRmR)a5R
SwRR:FRk0#_08DHFoOR;
RRRRRRRRQ:jRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;
0N0skHL0#CR$LM_D	NO_GLFRRFVp4zaRB:RFFlbM0CMRRH#0Csk;0
N0LsHkR0CGlO_NFbRVzRpa:4RRlOFbCFMMH0R#DR"k;0"
-S
-------------------------apz.-R--------------------------
--Bumvmhh azRpa
.RRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"Rj"2R;
RuRRmR)a5R
RRwSRRF:Rk#0R0D8_FOoH;R
RRQSRjRR:H#MR0D8_FOoH;R
RRQSR4RR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVp.zaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRa.:FROlMbFCRM0H"#RD"k0;-
-------------------------pdza-----------------------------B-
mmvuha hRapzdRR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjRj"2R;
RuRRmR)a5R
RRwSRRF:Rk#0R0D8_FOoH;R
RRQSRjRR:H#MR0D8_FOoH;R
RRQSR4RR:H#MR0D8_FOoH;R
RRQSR.RR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRad:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:dRRlOFbCFMMH0R#DR"k;0"
------------------------p--zRac-----------------------------m
Bvhum RhapczaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"j"jjR
2;RRRRuam)RR5
RRRSwRR:FRk0#_08DHFoOR;
RRRSQ:jRRRHM#_08DHFoOR;
RRRSQ:4RRRHM#_08DHFoOR;
RRRSQ:.RRRHM#_08DHFoOR;
RRRSQ:dRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVpczaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRac:FROlMbFCRM0H"#RD"k0;-
-------------------------p6zaR----------------------------B-
mmvuha hRapz6RR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjj";R2
RRRR)uma
R5RSRRR:wRR0FkR8#0_oDFH
O;RSRRRRQj:MRHR8#0_oDFH
O;RSRRRRQ4:MRHR8#0_oDFH
O;RSRRRRQ.:MRHR8#0_oDFH
O;RSRRRRQd:MRHR8#0_oDFH
O;RSRRRRQc:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRapz6RR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVp6zaRO:RFFlbM0CMRRH#"0Dk"-;
-------------------------apzn-R--------------------------
--
vBmu mhhpaRzRan
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjRj"2R;
RuRRmR)a5R
RRwSRRF:Rk#0R0D8_FOoH;R
RRQSRjRR:H#MR0D8_FOoH;R
RRQSR4RR:H#MR0D8_FOoH;R
RRQSR.RR:H#MR0D8_FOoH;R
RRQSRdRR:H#MR0D8_FOoH;R
RRQSRcRR:H#MR0D8_FOoH;R
RRQSR6RR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRan:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:nRRlOFbCFMMH0R#DR"k;0"
------------------------p--zRa(-----------------------------B

mmvuha hRapz(RR
RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj";R2
RRRR)uma
R5RSRRR:wRR0FkR8#0_oDFH
O;RSRRRRQj:MRHR8#0_oDFH
O;RSRRRRQ4:MRHR8#0_oDFH
O;RSRRRRQ.:MRHR8#0_oDFH
O;RSRRRRQd:MRHR8#0_oDFH
O;RSRRRRQc:MRHR8#0_oDFH
O;RRRRS6RQRH:RM0R#8F_Do;HO
RRRSnRQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:(RRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapz(RR:ObFlFMMC0#RHRk"D0
";-------------------------z-pa-UR----------------------------
m
Bvhum RhapUzaRR
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR
2;RRRRuam)RR5
RRRSwRR:FRk0#_08DHFoOR;
RRRSQ:jRRRHM#_08DHFoOR;
RRRSQ:4RRRHM#_08DHFoOR;
RRRSQ:.RRRHM#_08DHFoOR;
RRRSQ:dRRRHM#_08DHFoOR;
RRRSQ:cRRRHM#_08DHFoOR;
RRRSQ:6RRRHM#_08DHFoOR;
RRRSQ:nRRRHM#_08DHFoOR;
RRRSQ:(RRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVpUzaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRaU:FROlMbFCRM0H"#RD"k0;-
-------------------------v.zX-----------------------------
-
Bumvmhh azRvX
.RRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zXRB:RFFlbM0CMRRH#0Csk;-
-------------------------v.zX_apz6----------------------------
--
vBmu mhhvaRz_X.p6zaRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRa6:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.pnza-----------------------------
-
Bumvmhh azRvXp._zRan
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_pa:nRRlBFbCFMMH0R#sR0k
C;-------------------------z-vXp._z-a(-----------------------------B

mmvuha hRXvz.z_pa
(RRRRRuam)RS5
RRQj:MRHR8#0_oDFH
O;S4RQRH:RM0R#8F_Do;HO
1SRjRR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apz(RR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvz.z_pa-U-----------------------------
m
Bvhum Rhav.zX_apzURR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;SjR1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.pUzaRB:RFFlbM0CMRRH#0Csk;-
-------------------------v.zX_XvzU----------------------------
--
vBmu mhhvaRz_X.vUzXRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXv._zRXU:FRBlMbFCRM0H0#Rs;kC
------------------------v--z_X.v4zXn----------------------------
--
vBmu mhhvaRz_X.v4zXnRR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;SjR1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.v4zXnRR:BbFlFMMC0#RHRk0sC-;
-------------------------Xvz.z_vX-d.-----------------------------B

mmvuha hRXvz.z_vXRd.
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
S1:jRRRHM#_08DHFoOS;
R:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_vXRd.:FRBlMbFCRM0H0#Rs;kC
------------------------v--z-Xc-----------------------------B

mmvuha hRXvzcRR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;S.RQRH:RM0R#8F_Do;HORR
SQ:dRRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;S4R1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzRXc:FRBlMbFCRM0H0#Rs;kC
------------------------v--z-XU-----------------------------B

mmvuha hRXvzURR
RuRRmR)a5R
SQ:jRRRHM#_08DHFoOS;
RRQ4:MRHR8#0_oDFH
O;S.RQRH:RM0R#8F_Do;HORR
SQ:dRRRHM#_08DHFoOS;
RRQc:MRHR8#0_oDFH
O;S6RQRH:RM0R#8F_Do;HO
QSRnRR:H#MR0D8_FOoH;R
SQ:(RRRHM#_08DHFoOS;
RR1j:MRHR8#0_oDFH
O;S4R1RH:RM0R#8F_Do;HO
1SR.RR:H#MR0D8_FOoH;R
SmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvUzXRB:RFFlbM0CMRRH#0Csk;-
-------------------------v4zXn----------------------------
-
Bumvmhh azRvXR4nRR
RRmRu)5aR
QSRjRR:H#MR0D8_FOoH;R
SQ:4RRRHM#_08DHFoOS;
RRQ.:MRHR8#0_oDFHRO;
QSRdRR:H#MR0D8_FOoH;R
SQ:cRRRHM#_08DHFoOS;
RRQ6:MRHR8#0_oDFH
O;SnRQRH:RM0R#8F_Do;HO
QSR(RR:H#MR0D8_FOoH;R
SQ:URRRHM#_08DHFoOS;
RRQg:MRHR8#0_oDFH
O;S4RQjRR:H#MR0D8_FOoH;R
SQR44:MRHR8#0_oDFH
O;S4RQ.RR:H#MR0D8_FOoH;R
SQR4d:MRHR8#0_oDFH
O;S4RQcRR:H#MR0D8_FOoH;R
SQR46:MRHR8#0_oDFH
O;SjR1RH:RM0R#8F_Do;HO
1SR4RR:H#MR0D8_FOoH;R
S1:.RRRHM#_08DHFoOS;
RR1d:MRHR8#0_oDFH
O;SRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXR4n:FRBlMbFCRM0H0#Rs;kC
------------------------v--z.Xd-----------------------------B

mmvuha hRXvzdR.R
RRRR)uma
R5SjRQRH:RM0R#8F_Do;HO
QSR4RR:H#MR0D8_FOoH;R
SQ:.RRRHM#_08DHFoO
;RSdRQRH:RM0R#8F_Do;HO
QSRcRR:H#MR0D8_FOoH;R
SQ:6RRRHM#_08DHFoOS;
RRQn:MRHR8#0_oDFH
O;S(RQRH:RM0R#8F_Do;HO
QSRURR:H#MR0D8_FOoH;R
SQ:gRRRHM#_08DHFoOS;
RjQ4RH:RM0R#8F_Do;HO
QSR4:4RRRHM#_08DHFoOS;
R.Q4RH:RM0R#8F_Do;HO
QSR4:dRRRHM#_08DHFoOS;
RcQ4RH:RM0R#8F_Do;HO
QSR4:6RRRHM#_08DHFoOS;
RnQ4RH:RM0R#8F_Do;HO
QSR4:(RRRHM#_08DHFoOS;
RUQ4RH:RM0R#8F_Do;HO
QSR4:gRRRHM#_08DHFoOS;
RjQ.RH:RM0R#8F_Do;HO
QSR.:4RRRHM#_08DHFoOS;
R.Q.RH:RM0R#8F_Do;HO
QSR.Rd:RRHM#_08DHFoOS;
RcQ.RH:RM0R#8F_Do;HO
QSR.:6RRRHM#_08DHFoOS;
RnQ.RH:RM0R#8F_Do;HO
QSR.:(RRRHM#_08DHFoOS;
RUQ.RH:RM0R#8F_Do;HO
QSR.:gRRRHM#_08DHFoOS;
RjQdRH:RM0R#8F_Do;HO
QSRd:4RRRHM#_08DHFoO
;RSjR1RH:RM0R#8F_Do;HO
1SR4RR:H#MR0D8_FOoH;R
S1:.RRRHM#_08DHFoOS;
RR1d:MRHR8#0_oDFH
O;ScR1RH:RM0R#8F_Do;HO
mSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz.XdRB:RFFlbM0CMRRH#0Csk;-
-------------------------q-pz-----------------------------
-
Bumvmhh apRqzRR
RtRR )h Q5BRRRR
RRRRRRRRqR77:hRQa  t)=R:R;jR
RRRRRRRSzR1ARR:Q hatR ):4=RRR;
RRRRRRRRq177z:ARRaQh )t RR:=.
R;RRRRRSRRRRh :hRQa  t)=R:R;dR
RRRRRRRS RtRQ:Rhta  :)R=RRc;R
Sp: RRaQh )t RR:=6R;
RRRRRRRSBRzu:hRQa  t)=R:R;nR
RRRRRRRR7RBhRR:Q hatR ):(=RRR;
RRRRRRRRBBzu7:hRRaQh )t RR:=US;
RpvzaRR:Q hatR ):g=R;R
Sq_pzv m7RQ:Rhta  :)R=
RjRRRR2
;SRRRRuam)RS5
Rv1zRm:Rz#aR0D8_FOoH;R
SBamzRm:Rz#aR0D8_FOoH;SS
RRQj:hRQR8#0_oDFH
O;S4RQ:hRQR8#0_oDFH
O;SdRQ:hRQR8#0_oDFH
O;SQRBhQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFqVRp:zRRlBFbCFMMH0R#sR0k
C;----------------------------7Rww-----------------------------
-
Bumvmhh awR7wRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj;'2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rww:FRBlMbFCRM0H0#Rs;kC
---------------------------7 wwR--------------------------------
-
Bumvmhh awR7w
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSR RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRw :FRBlMbFCRM0H0#Rs;kC
------------------------w-7w-1R--------------------------------
m
Bvhum Rha71wwRR
RR RthQ )BRR5QahQ:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S1R a:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w1RR:BbFlFMMC0#RHRk0sC-;
-------------------------7--w w1-------------------------------------
-
Bumvmhh awR7wR1 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S1R a:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w1: RRlBFbCFMMH0R#sR0k
C;------------------------7)wwR--------------------------------
--
vBmu mhh7aRwRw)
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S)  1aRR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRw):FRBlMbFCRM0H0#Rs;kC
---------------------------7)ww -R----------------------------------
--
vBmu mhh7aRw w)RR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R1)  :aRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7)ww RR:BbFlFMMC0#RHRk0sC-;
-------------------------7--w-wu-------------------------------------
-
Bumvmhh awR7w
uRRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:uRRlBFbCFMMH0R#sR0k
C;-------------------------w-7wRu ---------------------------------------------B

mmvuha hRw7wu
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw wuRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--wRwB--------------------------------
m
Bvhum Rha7BwwRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R Bpq:)RRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7BwwRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--w wBR-------------------------------------------
m
Bvhum Rha7Bww RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wB: RRlBFbCFMMH0R#sR0k
C;-------------------------w-7w-hR-----------------------------B

mmvuha hRw7whRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj;'2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoO
;SSpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hwwRB:RFFlbM0CMRRH#0Csk;-
-----------------7hww -R------------------------------
--
vBmu mhh7aRw whRR
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
RRB :hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh: RRlBFbCFMMH0R#sR0k
C;-------------------------w7wh-1R--------------------------------
m
Bvhum Rha7hww1RR
RtRR )h Q5BRRQQhaL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
Ra1 RQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRh1:FRBlMbFCRM0H0#Rs;kC
----------------------------w7wh-1 -------------------------------------B

mmvuha hRw7whR1 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
S1R a:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
BSRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whR1 :FRBlMbFCRM0H0#Rs;kC
----------------------------w-7w-h)---------------------------------B

mmvuha hRw7wh
)RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
)SR a1 RQ:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRh):FRBlMbFCRM0H0#Rs;kC
---------------------------7hww)- R------------------------------------
m
Bvhum Rha7hww)
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
)SR a1 RQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
SBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w h)RB:RFFlbM0CMRRH#0Csk;-
--------------------------w-7w-hu-------------------------------------
-
Bumvmhh awR7wRhu
RRRRht  B)QRQ5RhRQa:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
Su1)  Ra:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwuwhRB:RFFlbM0CMRRH#0Csk;-
-------------------------7hwwu- R--------------------------------------------
m
Bvhum Rha7hwwu
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
uSR)  1aRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwuwh RR:BbFlFMMC0#RHRk0sC-;
----------------------------7hwwB-R------------------------------------------
-
Bumvmhh awR7wRhB
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwBwhRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--wBwh -R------------------------------------------B

mmvuha hRw7whRB 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH;SS
RiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRwBwh RR:BbFlFMMC0#RHRk0sC-;
-----------------------------7--p-R-----------------------------------------
m
Bvhum Rha7
pRRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7:pRRlBFbCFMMH0R#sR0k
C;------------------------- 7p---------------------------------
--
vBmu mhh7aRp
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rp :FRBlMbFCRM0H0#Rs;kC
----------------------------p-7B-R----------------------------------
-
Bumvmhh apR7BRR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB Rq):hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:BRRlBFbCFMMH0R#sR0k
C;-----------------------------B7p -R----------------------------------
-
Bumvmhh apR7B
 RRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HO
BSRp) qRQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH;R
SBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7 pBRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--p-uR---------------------------------
--
vBmu mhh7aRp
uRRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRR#:R0D8_FOoH;R
Su1)  :aRRRQh#_08DHFoO
;SS:RtRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu7pRB:RFFlbM0CMRRH#0Csk;-
--------------------------7--pRu ------------------------------------
m
Bvhum Rha7 puRR
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR
RRmRu)5aR
TSRRm:Rz#aR0D8_FOoH;SS
R:7RRRQh#_08DHFoOS;
R u)1R a:hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do;HO
BSR Q:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRu :FRBlMbFCRM0H0#Rs;kC
------------------------h7pR----------------------------------------
--
vBmu mhh7aRp
hRRRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRRQ:Rh0R#8F_Do;HOSR
StRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rph:FRBlMbFCRM0H0#Rs;kC
----------------------------p-7h- ----------------------------------B

mmvuha hRh7p RR
RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;RS
RuRRmR)a5R
STRR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHSO;
tSRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRh :FRBlMbFCRM0H0#Rs;kC
----------------------------p-7h-BR---------------------------------
--
vBmu mhh7aRpRhB
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7pBRR:BbFlFMMC0#RHRk0sC-;
----------------------------7Bph -R----------------------------------
-
Bumvmhh apR7hRB 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SBqp )RR:Q#hR0D8_FOoH;SS
R:tRRRQh#_08DHFoOS;
R:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7pB: RRlBFbCFMMH0R#sR0k
C;-----------------------------h7pu-R----------------------------------
-
Bumvmhh apR7h
uRRRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;SRRRRuam)RS5
R:TRRamzR8#0_oDFHSO;
7SRR#:R0D8_FOoH;R
Su1)  :aRRRQh#_08DHFoO
;SS:RtRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7puRR:BbFlFMMC0#RHRk0sC-;
----------------------------7uph -R----------------------------------
-
Bumvmhh apR7hRu 
RRRRht  B)QRQ5RhRQa:HRL0=R:R''4RS2;
RRRR)uma
R5SRRT:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
Su1)  :aRRRQh#_08DHFoO
;SSRRt:hRQR8#0_oDFH
O;S RB:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7hRu :FRBlMbFCRM0H0#Rs;kC
--------------------Q--A-zw------------------------------------
m
Bvhum RhaQwAzRR
RRmRu)5aR
RRRRmSRRm:Rz#aR0D8_FOoH;R
RRRRSQRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRARzw:FRBlMbFCRM0H0#Rs;kC
----------------------------m--A-zw-------------------------------------
-
Bumvmhh aARmz
wRRRRRuam)RR5
RSRRR:mRRamzR8#0_oDFH
O;RRRRSRRQ:hRQR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzmAwRR:BbFlFMMC0#RHRk0sC-;
---------------------------------a--A-zw-------------------------
-
Bumvmhh aARaz
wRRRRRuam)RR5
RSRRR:mRRamzR8#0_oDFH
O;RRRRSRRQ:hRQR8#0_oDFH
O;RRRRS RmhRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFaVRARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVawAzRB:RFFlbM0CMRRH#";m"
-
--------------------------m-QA-zw-----------------------------
--
vBmu mhhQaRmwAz
RRRR)uma
R5RRRRSRmR:zRmaRRR#_08DHFoOR;
RSRRQ:mRRmQhz#aR0D8_FOoH;R
RRSRRQ:RRRRQhR#RR0D8_FOoH;R
SRmRR :hRRRQhR#RR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRmwAzRB:RFFlbM0CMRRH#0Csk;-
------------------------------Q--7-7)-------------------------B

mmvuha hR7Q7)RR
RtRR )h Q5BR
jST_QQhaRR:LRH0:'=Rj
';S_T4QahQRL:RH:0R=jR''R
RR;R2SR
RRmRu)5aR
TSRjRR:mRza#_08DHFoOS;
RRT4:zRma0R#8F_Do;HOSR
S7RR:Q#hR0D8_FOoH;R
SB:piRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7Q7)RR:BbFlFMMC0#RHRk0sC
;
---------------------------------7Q7)-B--------------------------B

mmvuha hR7Q7)
BRRRRRt  h)RQB5SR
TQj_hRQa:HRL0=R:R''j;T
S4h_QQ:aRR0LHRR:='
j'RRRR2
;SRRRRuam)RS5
RRTj:zRma0R#8F_Do;HO
TSR4RR:mRza#_08DHFoO
;SSRR7:hRQR8#0_oDFH
O;SpRB :q)RRQh#_08DHFoO
;SSpRBiQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7B7)RB:RFFlbM0CMRRH#0Csk;-

-------------------------Q--7_7)v- v---------------------------------
--
vBmu mhhQaR7_7)vR v
 SthQ )B
R5S1St)R h:0R#soHMRR:="DVN#;C"
pSS1h) RRR:#H0sM:oR=0R"s"kC
;S2
mSu)5aR
TSSjRR:FRk0#_08DHFoO
;SS4STRF:Rk#0R0D8_FOoH;SS
S:7RRRHM#_08DHFoOS;
SpQBiRR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
WSSq)77RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SRRRS7)q7:)RRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ)77_vv RB:RFFlbM0CMRRH#0Csk;-

-----------------------------7-m7-)---------------------
vBmu mhhmaR7R7)
RRRRht  B)QR
5RRRRRRRRRapXBim_upRR:LRH0:'=RjR';-j-''H:)#oHMRoC8CkRF00bk;4R''N:wDMDHo8RCoFCRkk0b0RRRRRRRRR
RRRRRRmRBhq1ahQaRhRQa:0R#8F_DoRHO:'=Rj
'RRRRR2
;SRRRRuam)R
5RSRRRRRTj:zRma0R#8F_Do;HOSR
SRTRR4RR:mRza#_08DHFoO
;SSRRRRR7j:hRQR8#0_oDFH
O;SRRRRR74:hRQR8#0_oDFH
O;SRRRRRaX:hRQR8#0_oDFH
O;SRRRRiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR7R7):FRBlMbFCRM0H0#Rs;kC
-
------------------------------7m7)-B---------------------
m
Bvhum Rham)77BRR
RtRR )h Q5BRRR
RRRRRRXRaB_piuRmp:HRL0=R:R''j;-R-':j')HH#MCoR8RoCFbk0kR0;':4'wDNDHRMoCC8oR0Fkb
k0RRRRRRRRB1mhaaqhRQQhaRR:#_08DHFoO=R:R''j
RRRR
2;RRRRuam)RS5
RRRRT:jRRamzR8#0_oDFH
O;SRRRRRT4:zRma0R#8F_Do;HO
RSRRjR7RQ:Rh0R#8F_Do;HO
RSRR4R7RQ:Rh0R#8F_Do;HO
RSRRXRaRQ:Rh0R#8F_Do;HO
RSRRpRBiRR:Q#hR0D8_FOoH;R
SRBRRp) qRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR7B7)RB:RFFlbM0CMRRH#0Csk;-

-------------------------m--7_7)v- v---------------------------------
--Bumvmhh a7Rm7v)_ 
vRRRRRt  h)5QB
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)h:RRRs#0HRMo:"=R0Csk"R;
RRRRRaRRXiBp_pumRL:RH:0R=jR''-;R-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bk
RRRRRRRRpaBim_1z )BR#:R0MsHo=R:RT"71
W"RRRR2R;
RuRRmR)a5S
SRRTj:kRF00R#8F_Do;HOSS
SRRT4:kRF00R#8F_Do;HOSS
SRpaBiRR:H#MR0D8_FOoH;S
SRpuBiRR:H#MR0D8_FOoH;S
SR1)  :aRRRHM#_08DHFoOS;
SjR7RH:RM0R#8F_Do;HO
RSS7:4RRRHM#_08DHFoOS;
SXRaRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7v)_ :vRRlBFbCFMMH0R#sR0k
C;----------------------------------------- Q71-c------------------------------B

mmvuha hR Q71
cRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"S
2;S)uma
R5SRS7:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;S S)1R a:hRQR8#0_oDFH
O;SBSwp:iRRRQh#_08DHFoOS;
SpuBiRR:Q#hR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH;S
ST:.RRamzR8#0_oDFH
O;SdSTRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 cRR:BbFlFMMC0#RHRk0sC-;
------------------------- Q71vc_ -v---------------------------------
m
Bvhum RhaQ17 c _vvSR
oCCMs5HO
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)h:RRRs#0HRMo:"=R0Csk"2
S;u
Sm5)a
7SS,1)  :aRRRQh#_08DHFoOS;
SpBqQ:ARRRQh#_08DHFoOS;
SpQBiB,wpui,BRpi:hRQR8#0_oDFH
O;SqSW7R7):hRQR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
S7)q7:)RRRQh#_08DHFoOC_POs0F58.RF0IMF2Rj;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH;S
ST:.RRamzR8#0_oDFH
O;SdSTRm:Rz#aR0D8_FOoH
2SR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71vc_ :vRRlBFbCFMMH0R#sR0k
C;------------------------------------Q7eQ -m------------------------------B

mmvuha hRQQe7R m
RRRRht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7RR:Q#hR0D8_FOoH;S
S)  1aRR:Q#hR0D8_FOoH;S
SBQqpARR:Q#hR0D8_FOoH;S
SwiBpRQ:Rh0R#8F_Do;HO
uSSBRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRe Q7mRR:BbFlFMMC0#RHRk0sC-;
---------------------------------7-Q -1U------------------------------------
m
Bvhum RhaQ17 URR
RtRR )h Q5BR
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
pSS1h) RRR:#H0sM:oR=0R"s"kC
RRRR
2;RRRRuam)RS5
S)7, a1 RQ:Rh0R#8F_Do;HO
BSSqApQRQ:Rh0R#8F_Do;HO
wSSB,piuiBpRQ:Rh0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do;HO
TSS.RR:mRza#_08DHFoOS;
SRTd:zRma0R#8F_Do;HO
TSScRR:mRza#_08DHFoOS;
SRT6:zRma0R#8F_Do;HO
TSSnRR:mRza#_08DHFoOS;
SRT(:zRma0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ R1U:FRBlMbFCRM0H0#Rs;kC
------------------------7-Q _1Uv- v-------------------------
--
vBmu mhhQaR7U 1_vv RR
RR RthQ )B
R5SRRRR)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7 ,)1R a:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;SBSwpQi,B,piuiBpRQ:Rh0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do;HO
TSS.RR:mRza#_08DHFoOS;
SRTd:zRma0R#8F_Do;HO
TSScRR:mRza#_08DHFoOS;
SRT6:zRma0R#8F_Do;HO
TSSnRR:mRza#_08DHFoOS;
SRT(:zRma0R#8F_Do;HO
WSSq)77RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SqS)7R7):MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 U _vvRR:BbFlFMMC0#RHRk0sC-;
------------------------------------- Q71-4j---------------------------------B

mmvuha hR Q71R4j
RRRRht  B)QRS5
RRRRt 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 RhR:0R#soHMRR:="k0sCR"
R2RR;R
RRmRu)5aR
7SS,1)  :aRRRQh#_08DHFoOS;
SpBqQ:ARRRQh#_08DHFoOS;
SpwBiB,up:iRRRQh#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoOS;
SRT.:zRma0R#8F_Do;HO
TSSdRR:mRza#_08DHFoOS;
SRTc:zRma0R#8F_Do;HO
TSS6RR:mRza#_08DHFoOS;
SRTn:zRma0R#8F_Do;HO
TSS(RR:mRza#_08DHFoOS;
SRTU:zRma0R#8F_Do;HO
TSSgRR:mRza#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 4:jRRlBFbCFMMH0R#sR0k
C;------------------------- m1)-c-----------------------------
m
Bvhum Rham)1 cSR
t  h)RQB5S
St 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 :hRRs#0HRMo:"=R0Csk"R;
RRRRR]RRW:pRRs#0HRMo:"=RV#NDCR";-0-"s"kC;VR"NCD#"R
RRRRRRXRaB_piuRmp:HRL0=R:R''jR'--j)':HM#Ho8RCoFCRkk0b0';R4w':NHDDMCoR8RoCFbk0kS0
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SjaXRH:RM0R#8F_Do;HO
aSSX:4RRRHM#_08DHFoOS;
SpuBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SwiBpRH:RM0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR1c )RB:RFFlbM0CMRRH#0Csk;-
--------------m--1c )_vv --------------------------------
m
Bvhum Rham)1 c _vvSR
t  h)RQB5S
St 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 :hRRs#0HRMo:"=R0Csk"S;
Sp]WR#:R0MsHo=R:RN"VD"#C;R
RRRRRRXRaB_piuRmp:HRL0=R:R''j;'--j)':HM#Ho8RCoFCRkk0b0';R4w':NHDDMCoR8RoCFbk0kR0
RRRRRaRRB_pi1)mzB: RRs#0HRMo:"=R7WT1"2
S;u
SmR)a5S
S7:jRRRHM#_08DHFoOS;
SR74:MRHR8#0_oDFH
O;S.S7RH:RM0R#8F_Do;HO
7SSdRR:H#MR0D8_FOoH;S
SaRXj:MRHR8#0_oDFH
O;SXSa4RR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SBSap:iRRRHM#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1)vc_ :vRRlBFbCFMMH0R#sR0k
C;--------------------m7eQ -m---------------------------------
m
Bvhum Rham7eQ 
mRSht  B)Q5S
St 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 :hRRs#0HRMo:"=R0Csk"2
S;u
SmR)a5S
S7:jRRRHM#_08DHFoOS;
SR74:MRHR8#0_oDFH
O;S.S7RH:RM0R#8F_Do;HO
7SSdRR:H#MR0D8_FOoH;S
S7:cRRRHM#_08DHFoOS;
SR76:MRHR8#0_oDFH
O;SnS7RH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSwp:iRRRHM#_08DHFoOS;
S:TRRamzR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVeRmQm7 RB:RFFlbM0CMRRH#0Csk;-
------------------1-m -)U---------------------------------
-
Bumvmhh a1Rm R)U
RRRRht  B)QRR5
RSRRt 1)hRR:#H0sM:oR=VR"NCD#"R;
RSRRp 1)hRR:#H0sM:oR=0R"s"kC;R
RRRRRRWR]pRR:#H0sM:oR=VR"NCD#"R;
RRRRRaRRXiBp_pumRL:RH:0R=jR''-R-':j')HH#MCoR8RoCFbk0kR0;':4'wDNDHRMoCC8oR0FkbRk0RR
R2R;
RuRRmR)a5R
RRRRRRjS7RH:RM0R#8F_Do;HO
RRRRRRRSR74:MRHR8#0_oDFH
O;RRRRRSRR7:.RRRHM#_08DHFoOR;
RRRRR7RSdRR:H#MR0D8_FOoH;R
RRRRRRcS7RH:RM0R#8F_Do;HO
RRRRSRR7:6RRRHM#_08DHFoOR;
RRRRR7RSnRR:H#MR0D8_FOoH;R
RRRRRR(S7RH:RM0R#8F_Do;HO
RRRRRRRSjaXRH:RM0R#8F_Do;HO
RRRRXSa4RR:H#MR0D8_FOoH;R
SRaRRX:.RRRHM#_08DHFoOS;
RRRRaRXd:MRHR8#0_oDFH
O;SRRRRpuBiRR:H#MR0D8_FOoH;R
SR)RR a1 RH:RM0R#8F_Do;HO
RSRRBRwp:iRRRHM#_08DHFoOR;
RRRRRTRSjRR:mRza#_08DHFoOR;
RRRRRTRS4RR:mRza#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 URR:BbFlFMMC0#RHRk0sC-;
----------------m)1 U _vv--------------------------------B

mmvuha hR m1)vU_ 
vRSht  B)Q5S
St 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 :hRRs#0HRMo:"=R0Csk"S;
Sp]WR#:R0MsHo=R:RN"VD"#C;R
RRRRRRXRaB_piuRmp:HRL0=R:R''j;R
RRRRRRBRap1i_mBz) RR:#H0sM:oR=7R"T"1W
;S2
mSu)5aR
7SSjRR:H#MR0D8_FOoH;S
S7:4RRRHM#_08DHFoOS;
SR7.:MRHR8#0_oDFH
O;SdS7RH:RM0R#8F_Do;HO
7SScRR:H#MR0D8_FOoH;S
S7:6RRRHM#_08DHFoOS;
SR7n:MRHR8#0_oDFH
O;S(S7RH:RM0R#8F_Do;HO
aSSX:jRRRHM#_08DHFoOS;
S4aXRH:RM0R#8F_Do;HO
aSSX:.RRRHM#_08DHFoOS;
SdaXRH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSwp:iRRRHM#_08DHFoOS;
SpaBiRR:H#MR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 U _vvRR:BbFlFMMC0#RHRk0sC-;
-----------------m--14 )j-----------------------------------
m
Bvhum Rham)1 4
jRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sCS"
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SR7c:MRHR8#0_oDFH
O;S6S7RH:RM0R#8F_Do;HO
7SSnRR:H#MR0D8_FOoH;S
S7:(RRRHM#_08DHFoOS;
SR7U:MRHR8#0_oDFH
O;SgS7RH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SBSwp:iRRRHM#_08DHFoOS;
S:TRRamzR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rm j)4RB:RFFlbM0CMRRH#0Csk;-
------------------m-Q7q pY-----------------------------------
m
Bvhum RhaQ m7pRqY
 SthQ )BRR5R1B_aQqaBp_7YRR:HCM0oRCs:j=R2-;R-~Rj4
.(S)uma
R5SQS7RQ:Rh0R#8F_Do;HO
1SS7uaqRQ:Rh0R#8F_Do;HO
1SS Rah:hRQR8#0_oDFH
O;SqSepRz :hRQR8#0_oDFH
O;SmS7Rm:Rz#aR0D8_FOoH;S
S7:wRRamzR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVmRQ7q pYRR:BbFlFMMC0#RHRk0sC-;
-----------------Q-- -v---------------------------------
m
Bvhum RhaQR v
 SthQ )BS5
ShWQ1 QZR#:R0MsHo=R:Rv"1q"pp;S
St 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 RhR:0R#soHMRR:="k0sCS"
2S;
uam)RS5
S:7RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
vSSB:piRRHM#_08DHFoOS;
StpqRF:Rk#0R0D8_FOoH;S
Sp7 qRF:Rk#0R0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQR v:FRBlMbFCRM0H0#Rs;kC
-----------------------)-mv-------------------------
--
vBmu mhh)aRm
vRRRRRt  h)RQB5SR
RaAQ_7WQa:]RR0HMCsoCR4:=;SS
Rq) 7m_v7: RR0LHRR:=';j'
RRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRRRRR
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsj.,d2S;
RiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoOR;
RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
Sq:7RRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)Rmv:FRBlMbFCRM0H0#Rs;kC
----------------------------)--mgvXR--------------------------------------------
-
Bumvmhh amR)vRXg
RRRRht  B)QR
5RRRRRA_QaWaQ7]RR:HCM0oRCs:;=g
RRRRq) 7m_v7: RR0LHR':=j
';RRRRA_pi1R p:HRL0C_POs0FRR:="jjj"R;
R)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBRRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
R
RRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
BSRpRi,Bm ,B) , a1 , W)RH:RM0R#8F_Do;HO
RRRRASRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
qSR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRmgvXRB:RFFlbM0CMRRH#0Csk;-

-----------------u-1-------------------------------------
--Bumvmhh auR1RR
RR RthQ )B
R5SQRAaQ_W7Ra]:MRH0CCos=R:dR.;-4-R,,R.RRc,U4,Rnd,R.R
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)RWQ_a v m7RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiB,R B,m  ,)1, aWR) :MRHR8#0_oDFH
O;S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds54FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR1RB:RFFlbM0CMRRH#0Csk;-

-------------------------1--u-Xg-------------------------------------
-
Bumvmhh auR1X
gRRRRRt  h)RQB5SR
RaAQ_7WQa:]RR0HMCsoCRg:=;R
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)RWQ_a v m7RL:RHP0_CFO0s=R:""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRR
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoOS;
RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2
RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR1X:gRRlBFbCFMMH0R#sR0k
C;



---------------------------------7-1u-A--------------------------------------m
Bvhum Rha1A7uRR
RR RthQ )BRR5
RSRRQRAaQ_W7_a]jRR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.SRRRRaAQ_7WQa4]_RH:RMo0CC:sR=;4nRR--4.,R,,RcRRU,4Rn,dS.
RRRR)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CRRRRRRRRA_pi1_ pjRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRRiAp_p1 _:4RR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SRBRRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  RaA:MRHR8#0_oDFH
O;SRRRRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRRRRRiAp1q p,iAp1A pRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SRRRRR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu17ARR:BbFlFMMC0#RHRk0sC
;
---------------------------------7-1uAXg-------------------------------------
--Bumvmhh a7R1uAXgRR
RR RthQ )BRR5
RSRRQRAaQ_W7_a]jRR:HCM0oRCs:U=4;-R-RRg,4RU,dSn
RRRRA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4,nRd
RSRR R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SRARRp1i_ jp_RL:RHP0_CFO0s=R:Rj"jj
";SRRRRiAp_p1 _:4RR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
RRRRRR2R;
RuRRmR)a5R
SR7RRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SRRRRiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 ARR:H#MR0D8_FOoH;R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRRARRp i1pAq,p i1p:ARRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SR7RRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF1VR7guXARR:BbFlFMMC0#RHRk0sC
;
----------------------------7-uA-------------------------------------
-
Bumvmhh auR7ARR
RtRR )h Q5BR
RSSA_QaWaQ7]R_j:MRH0CCos=R:4Rn;
RSSA_QaWaQ7]R_4:MRH0CCos=R:4Rn;
RSS)7 q_7vm :jRR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
RSS)7 q_7vm :4RR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
RSSWa)Q m_v7R j:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RSSWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RRRRASRp1i_ jp_RL:RHP0_CFO0s=R:Rj"jj
";RRRRSpRAi _1pR_4:HRL0C_POs0FRR:="jjj"R;
RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSSQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
j"RRRR2R;
RuRRmR)a5S
SRq7m,A7mRF:Rk#0R0D8_FOoH_OPC05Fs486RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,42S;
SpRBiBq,p,iARqB ,AB , mBqB,m )A, a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRRRSA1pi ,pqA1pi RpA:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRu:ARRlBFbCFMMH0R#sR0k
C;
----------------------------X7ug-A--------------------------------------m
Bvhum Rha7guXARR
RtRR )h Q5BRRR
SRARRQWa_Q]7a_:jRR0HMCsoCR4:=U-;R-,RgR
4USRRRRaAQ_7WQa4]_RH:RMo0CC:sR=;4URR--g4,RUR
SR)RR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSRRRRq) 7m_v7R 4:HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SRWRR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CSRRRRQW)av _m47 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRRRRRpRAi _1pR_j:HRL0C_POs0FRR:="jjj"R;
RRRRRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
RRRR
2;RRRRuam)RS5
RRRR7,mq7RmA:kRF00R#8F_Do_HOP0COF4s5(FR8IFM0RRj2:O=RF_MP#_08DHFoOC_POs0F54j,U
2;SRRRRiBpqp,BiRA,B, qB, AmqB , mBA ,)1q a,1)  ,aAWq) , W)ARR:H#MR0D8_FOoH;R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
RRRR7RQq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;RRRRRRRRA1pi ,pqA1pi RpA:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RRRR7RQA:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRX7ug:ARRlBFbCFMMH0R#sR0k
C;







---------------------------------7-1u---------------------------------------
m
Bvhum Rha1R7u
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
S7:QRRRHM#_08DHFoOC_POs0F5Rd48MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV1R7u:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------1X7ug---------------------------------------
m
Bvhum Rha1X7ugRR
RtRR )h Q5BRRR
SA_QaWaQ7]R_j:MRH0CCos=R:4RU;-g-R,UR4,nRd
ASRQWa_Q]7a_:4RR0HMCsoCR4:=U-;R-,RgR,4UR
dnS R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SA_pi1R p:HRL0C_POs0FRR:="jjj"R;
RRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRRR
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRARRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
7SRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF1VR7guXRB:RFFlbM0CMRRH#0Csk;

S---------------------------------1-s7-u--------------------------------------m
Bvhum Rhasu17RR
RR RthQ )BRR5
ASRQWa_Q]7a_:jRR0HMCsoCR4:=n-;R-,R4RR.,cU,R,nR4,.Rd
ASRQWa_Q]7a_:4RR0HMCsoCR4:=n-;R-,R4RR.,cU,R,nR4,.Rd
)SR _q7v m7RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8RC
RRRRA_pi1R p:HRL0C_POs0FRR:="jjj"R;
RRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"R
RRRRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
BSRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  RaA:MRHR8#0_oDFH
O;S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRARRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
7SRQRR:H#MR0D8_FOoH_OPC05Fsd84RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR1R7u:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------su17X-g--------------------------------------m
Bvhum Rhasu17X
gRRRRRt  h)RQB5SR
RaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUd,RnR
SA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4,nRd
)SR _q7v m7RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
RiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1a:ARRRHM#_08DHFoOS;
Rqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rs7guXRB:RFFlbM0CMRRH#0Csk;



-
----------------------mb)v----------------------------m
Bvhum Rhabv)mRR
RR RthQ )BRR5
RSRRQRAaQ_W7Ra]:MRH0CCos=R:4
;SSRRRRq) 7m_v7: RR0LHRR:=';j'
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRRRR
RRRR
2;RRRRuam)RS5
RRRR7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
RSRRpRBiB,R m,RBR ,)  1aRR:H#MR0D8_FOoH;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFbVR)Rmv:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------bv)mX-gR--------------------------------------------
vBmu mhhbaR)XmvgRR
RtRR )h Q5BRRR
RRRRRRQRAaQ_W7Ra]:MRH0CCos=R:gR;
RRRRR)RR _q7v m7RL:RH:0R=''j;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hRB
RRRRRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRR

R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SpRBiB,R m,RBR ,)  1aRR:H#MR0D8_FOoH;R
Sq:7RRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVbv)mX:gRRlBFbCFMMH0R#sR0k
C;



---------------------s--)-mv-------------------------
--Bumvmhh a)Rsm
vRRRRRt  h)RQB5SR
RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SR
SR)RR _q7v m7RL:RH:0R=jR''R;
RRRRRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SRBRRpRi,BR ,m,B R1)  :aRRRHM#_08DHFoOR;
RSRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR)Rmv:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------sv)mX-gR--------------------------------------------
vBmu mhhsaR)XmvgRR
RtRR )h Q5BRRR
RRRRRRQRAaQ_W7Ra]:MRH0CCos=R:gR;
RRRRR)RR _q7v m7RL:RH:0R=''j;R
RRRRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
RRRRRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
R
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB,BRm ),R a1 RH:RM0R#8F_Do;HO
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV)RsmgvXRB:RFFlbM0CMRRH#0Csk;


----------------------------7-u--------------------------------------B

mmvuha hRR7u
RRRRht  B)QRS5
SQRAaQ_W7_a]jRR:HCM0oRCs:n=4;SR
SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;SR
S R)qv7_mj7 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S)RWQ_a v m7jRR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
S)RWQ_a v m74RR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8RC
RSRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBS
SRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj
RRRR
2;RRRRuam)RS5
SmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R468MFI0jFR2O:=F_MP#_08DHFoOC_POs0F54j,n
2;SBSRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;SqSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuRR:BbFlFMMC0#RHRk0sC
;
----------------------------7guX-------------------------------------
--
vBmu mhh7aRuRXg
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:U=4;-R-RRg,4SU
RaAQ_7WQa4]_RH:RMo0CC:sR=;4URR--g4,RUR
S)7 q_7vm :jRR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
)SR _q7v m74RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)RWQ_a v m7jRR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
RQW)av _m47 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RR
RRRRRR2R;
RuRRmR)a5R
S7,mq7RmA:kRF00R#8F_Do_HOP0COF4s5(FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,24U;R
SBqpi,iBpAB,R Bq, mA,B, qmAB ,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
Rq7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuRXg:FRBlMbFCRM0H0#Rs;kC
-
------------------------------q-)v14n4------------------------
--
vBmu mhh)aRqnv41
4RRRRRt  h)RQB5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj";R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S)SW RR:H#MR0D8_FOoH;S
Sq:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S7:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnR14:FRBlMbFCRM0H0#Rs;kC
--------------------------------v)q4.n1-------------------------
-
Bumvmhh aqR)v14n.RR
RtRR )h Q5BRRQQhaR_j:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
SRRRRRRRRRQQhaR_4:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jjRR
RRRRRRRRRR;R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
BSSp:iRRRHM#_08DHFoOS;
S W)RH:RM0R#8F_Do;HO
qSS7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
7SSQRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n.RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41-c-------------------------
m
Bvhum Rha)4qvnR1c
RRRRht  B)Q5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"S;
RRRRRRRRRQQhaR_4:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
SRRRRRRRRQahQ_:.RR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RRRRRRRRRRRRhRQQda_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R
RRRRRRRRRR
2;RRRRuam)RS5
SR7m:kRF00R#8F_Do_HOP0COFds5RI8FMR0FjR2;
BSSp:iRRRHM#_08DHFoOS;
S W)RH:RM0R#8F_Do;HO
qSS7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
7SSQRR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14ncRR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv4147u-------------------------R-
Rm
Bvhum Rha)4qvnu174RR
RtRR )h QRB5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jjRj"2R;
RuRRmR)a5S
S7:mRR0FkR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
SWR) :MRHR8#0_oDFH
O;SqSW7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
)SSq:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S7:QRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu174RR:BbFlFMMC0#RHRk0sC-;
-----------------------------)--qnv41.7u-------------------------
-
Bumvmhh aqR)v14n7Ru.
RRRRht  B)QRQ5Rh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";SRRRRRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjjR"
RRRRRRRRR2RR;R
RRmRu)5aR
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RSRRpRBiRR:H#MR0D8_FOoH;R
SRWRR): RRRHM#_08DHFoOS;
RRRRWRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
RRRR)Rq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
RRRR7:QRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRqnv41.7uRB:RFFlbM0CMRRH#0Csk;-
------------------------------q-)v14n7-uc-------------------------B

mmvuha hRv)q47n1u
cRRRRRt  h)RQB5hRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"S;
RRRRRRRRRhRQQ4a_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R;
RRRRRRRRRRRRRQQhaR_.:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
RRRRRRRRRRRRRQahQ_:dRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj
j"RRRRRRRRRRRR2R;
RuRRmR)a5S
S7:mRR0FkR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
S7WqRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;SqS)7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
7SSQRR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n7Ruc:FRBlMbFCRM0H0#Rs;kC
-
------------------------------m-)v-4n----------------------------
vBmu mhh)aRmnv4RR
RR RthQ )BRR5QahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jjRj"2R;
RuRRmR)a5S
RRRRR7:mRR0FkR8#0_oDFH
O;SRRRRRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4mvnRR:BbFlFMMC0#RHRk0sC
;
---------------------wAzt---------------------------
m
Bvhum RhaAtzwRR
Ruam)5R
RRmRSRF:Rk#0R0D8_FOoH;R
RRQRSRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRAw:tRRlBFbCFMMH0R#sR0k
C;-----------------wAz1--------------------B

mmvuha hRwAz1RR
RuRRmR)a5R
RRRRRRmRRRF:Rk#0R0D8_FOoH;R
RRRRRRQRRRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRAw:1RRlBFbCFMMH0R#sR0k
C;---------------------h-t7----------------
-
Bumvmhh ahRt7RR
RuRRmR)a5R
RRRRStRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVtRh7:FRBlMbFCRM0H0#Rs;kC
--------------------B-eB------------------------B

mmvuha hRBeBRR
RRmRu)5aR
RRRReSRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFeVRB:BRRlBFbCFMMH0R#sR0k
C;
----------------m--1-B--------------------------B-
mmvuha hRBm1RR
RR RthQ )B
R5RRRRRRRRwT) _e7QRH:RMo0CC:sR=jR4jR;R-~-.4,.UF$MDRCCPMkRMlR
RRRRRR R7e QBR#:R0MsHo=R:RW"t.4q-U-"R-.tWqU-4,.tWq6-6,.tWq4)-UR
RR;R2
RRRR)uma
R5SRRRRBm1mRza:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1RmBRR:BbFlFMMC0#RHRk0sCS;

----------------h-Qe--------------------------------
-
Bumvmhh ahRQeRR
RuRRmR)a5R
RRRRSmRR:mRza#_08DHFoOR;
RSRRR:QRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQRhe:FRBlMbFCRM0H0#Rs;kC
-
--------------7--p-p------------------------------
--Bumvmhh apR7pR
RR RthQ )BR5
RRRRR7RRpwp_m )BRH:RMo0CC:sR=;Rj-:-4RsVFODCRFRO	NRM8OCF8;:RjR8OFCF/DOo	RCsMCN80CRFVslpR7pFRDFRb
RRRRR7RRQ1e_ :pRR0LHRR:=';4'-,-jMlFsNDDRFRO	lCF8;,R4V0N#RODF	FRl8SC
RRRRB m71pBqR1:Rah)Qt=R:Rj"jj-";-4jjRjj4R4j4Rj4jR44jRj44R444
RRRRRRRRq1Bph_ R1:Rah)Qt=R:Rs"0k-C"-k0sCN,VD
#CRRRR2R;
RuRRm5)a
RRRRRRRRiBpQQh:h0R#8F_Do:HO=''j;R
RRRRRRaR1mRu:Q#MR0D8_FOoH:j=''R;
RRRRR)RR a1 RQ:RM0R#8F_Do:HO=''j;R
RRRRRRuRz7hhBa:pRRRQM#_08DHFoO':=j
';RRRRRRRRpimBRm:Rz#aR0D8_FOoH;R
RRRRRRaR1 :uRRamzR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R
RR2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRp7pRB:RFFlbM0CMRRH#0Csk;


-----------------eap7Q1_A-zw--------------------------------
m
Bvhum Rhaa7pe1A_QzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH;R
RRRRRRARQRQ:Rh0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFReap7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1A_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------eap7m1_A-zw--------------------------------
m
Bvhum Rhaa7pe1A_mzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRm:ARRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH
RRRRRRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpRae_71mwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFReap7m1_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------p-ae_71awAz---------------------------------B

mmvuha hReap7a1_A
zwRRRRuam)RR5
RSRRRRmR:zRmaRRR#_08DHFoOR;
RSRRRRmA:zRma0R#8F_Do;HO
RRRRRRSQ:RRRRQhR#RR0D8_FOoH;R
SRRRRmR h:hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGFaVRp1e7_zaAwRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpRae_71awAzRB:RFFlbM0CMRRH#"Rm,m;A"
-
--------------a--p1e7_AQmz-w------------------------------
--
vBmu mhhaaRp1e7_AQmzRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSQRmA:hRQmRza#_08DHFoOR;
RRRRRRRRQ:mRRmQhz#aR0D8_FOoH;R
RRSRRRRQR:hRQRRRR#_08DHFoOS;
RRRRRhm RQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVa7pe1m_QARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1m_QARzw:FRBlMbFCRM0H"#RQRm,Q"mA;-

---------------- 7pe1A_Qz-w------------------------------
--
vBmu mhh aRp1e7_zQAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do;HO
RRRRRRRRRQA:hRQR8#0_oDFHRO
RRRRR2RR;M
C8mRBvhum ;ha
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFV 7pe1A_Qz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMF VRp1e7_zQAwRR:BbFlFMMC0#RHR,"QR"QA;-

---------------- 7pe1A_mz-w------------------------------
--
vBmu mhh aRp1e7_zmAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRmRRARR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7m1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_mz:wRRlBFbCFMMH0R#mR",ARm"
;
-----------------e p7a1_A-zw--------------------------------
m
Bvhum Rha 7pe1A_azRw
RuRRmR)a5R
RRRRSm:RRRamzR#RR0D8_FOoH;R
RRRRSm:ARRamzR8#0_oDFH
O;RRRRRQSRRRR:QRhRR0R#8F_Do;HO
RSRRmRR :hRRRQhR#RR0D8_FOoH
RRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpR e_71awAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRe p7a1_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------p- e_71QzmAw--------------------------------
-
Bumvmhh apR e_71QzmAwR
RRmRu)5aR
RRRRmSRRRR:mRzaR0R#8F_Do;HO
RRRRQSRm:ARRmQhz#aR0D8_FOoH;R
RRRRRRQRRmRR:Qzhma0R#8F_Do;HO
RRRRRRSQ:RRRRQhR#RR0D8_FOoH;R
SRRRRmR h:hRQRRRR#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;RRRRNs00H0LkC$R#MD_LN_O	LRFGF VRp1e7_AQmz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMF VRp1e7_AQmz:wRRlBFbCFMMH0R#QR"mQ,Rm;A"
-
--------------------------q-u7U74-------------------------------------
--Bumvmhh aqRu7U74
oSSCsMCH
O5SRSRR)Rq :tRR0LHRR:=';j'-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SRRRRAt) RL:RH:0R=jR''
;RSRSRRmR1)R t:HRL0=R:R''j;S
SRRRRq_771RzA:HRL0=R:R''j;R
RRRRRRRRRRqRu7)7_ a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-Rh1YB1,qY
hBRRRRRRRRRRRRAp1 _7vm RR:LRH0:'=R4-'R-4R""#:RE0HV,jR""b:RNDsNDRCDHkMb03RA
RSRR;R2
RRRRRRR
RRRRRRRRsbF0S5
SRRRR:qRRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SRRRR:ARRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
SRRRR q1pRR:H#MR0D8_FOoH;S
SRRRRBB ,p)i, a1 RH:RM0R#8F_Do;HO
RSSR1RRQA,1QRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SRRRR11m,A:mRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0FjR2
RSRR2 ;
hB7Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqRu7U74RB:RFFlbM0CMRRH#0Csk;-

-------------------------u--qg77-------------------------------------
--Bumvmhh aqRu7
7gRRRRRRRRoCCMs5HO
RSSRqRR)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8SC
SRRRR A)tRR:LRH0:'=RjR';
RSSR1RRmt) RL:RH:0R=jR''S;
SRRRR7q7_A1zRL:RH:0R=jR''R;
RRRRRRRRRuRRq_77)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-YR1hqB,1BYh
RRRRRRRRRRRR A1pm_v7: RR0LHRR:='R4'-"-R4R":#VEH0",RjR":bNNsDDDCRbHMkA0R3R
SR2RR;R
RRRRRRRR
RSRRb0FsRS5
SRRRR:qRRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
SRRRRARR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
RSSRqRR1R p:MRHR8#0_oDFH
O;SRSRR RB,iBp,1)  :aRRRHM#_08DHFoOS;
SRRRR,1Q1RAQ:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SRRRR,1m1RAm:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;SRSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0sR5U8MFI0jFR2R
SR2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7uq7:gRRlBFbCFMMH0R#sR0k
C;
----------------------------pvzaggX-------------------------------------m
Bvhum Rhavazpg
XgSCSoMHCsOS5
SRRRR q)tRR:R0LHRR:=';j'RR--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CSRSRR)RA :tRRHRL0=R:R''j;S
SRRRRm_za)R t:LRRH:0R=jR''S;
SRRRRuuQ  _)tRR:R0LHRR:=';j'
RSSRqRR1hQt_t) RR:RLRH0:'=Rj
';SRSRR1RAQ_th)R t:LRRH:0R=jR''R;
RRRRRRRRR1RRm)q_ :tRRHRL0=R:R''j;SR
SRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
RRRR2
;
RRRRSsbF0
R5SRSRR,Rq1RQq:MRHR8#0_oDFHPO_CFO0sR5U8MFI0jFR2S;
SRRRR1A,Q:ARRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S
SRRRRqt1QhA,R1hQtRH:RM0R#8F_Do;HO
RRRRRRRRRRRR q1p1,A :pRRRHM#_08DHFoOS;
SRRRRRB :MRHR8#0_oDFH
O;SRSRRpRBiRR:H#MR0D8_FOoH;S
SRRRR)  1aRR:H#MR0D8_FOoH;S
SRRRR7amzRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj;R
RRRRRRRRRRmR1qm,1ARR:FRk0#_08DHFoOC_POs0F58URF0IMF2Rj
RSRR;R2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpgRXg:FRBlMbFCRM0H0#Rs;kC
-
--------------------------z-vpUa4X-4U-------------------------------------
-
Bumvmhh azRvpUa4X
4URRRRoCCMs5HO
qSS)R t:LRRH:0R=jR''-;R-'RRjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SAt) RR:RLRH0:'=Rj
';SzSma _)tRR:R0LHRR:=';j'
uSSQ_u )R t:LRRH:0R=jR''S;
SQq1t)h_ :tRRHRL0=R:R''j;S
SAt1Qh _)tRR:R0LHRR:=';j'
RRRRRRRRq1m_t) RR:RLRH0:'=Rj
';SzSvp)a_ a1 _7vm RR:#H0sM:oR=1R"Y"hBRR--1BYh,1RqY
hBS
2;
FSbs50R
qSS,q1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
ASS,A1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
qSS1hQt,1RAQRth:MRHR8#0_oDFH
O;RRRRRRRRqp1 , A1pRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
7SSmRza:kRF00R#8F_Do_HOP0COFds56FR8IFM0R;j2
RRRRRRRRq1m,A1mRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazp44UXURR:BbFlFMMC0#RHRk0sC
;
----------------------------vazpddnXn---------------------------------------
vBmu mhhvaRzdpannXd
CSoMHCsOS5
S q)tRR:R0LHRR:=';j'RR--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CS)SA :tRRHRL0=R:R''j;S
Smjza_t) RR:RLRH0:'=Rj
';SzSma)4_ :tRRHRL0=R:R''j;S
Su Qu_t) RR:RLRH0:'=Rj
';S1SqQ_th)R t:LRRH:0R=jR''S;
SQA1t)h_ :tRRHRL0=R:R''j;S
Svazp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-YR1hRB,qh1YB2
S;S

b0FsRS5
S:qRRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
S:ARRRHM#_08DHFoOC_POs0F5Rd68MFI0jFR2S;
SQq1tRh,At1QhRR:H#MR0D8_FOoH;S
SB: RRRHM#_08DHFoOS;
SiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
7SSmRza:kRF00R#8F_Do_HOP0COF(s54FR8IFM0R
j2S
2; Rh7Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRzdpannXdRB:RFFlbM0CMRRH#0Csk;-

-------------------------v--zqpapnzdX-4U-------------------------------------B-
mmvuha hRpvzazqpd4nXUo
SCsMCH
O5S)Sq :tRRHRL0=R:R''j;-R-RjR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
ASS)R t:LRRH:0R=jR''S;
S B)tRR:R0LHRR:=';j'
mSSz)a_ :tRRHRL0=R:R''j;S
Su Qu_t) RR:RLRH0:'=Rj
';S1SqQ_th)R t:LRRH:0R=jR''S;
SQA1t)h_ :tRRHRL0=R:R''j;R
RRRRRRBRqBqpm7 _)t:jRR0LHRR:=';j'
RRRRRRRRBqBp7mq_t) 4RR:LRH0:'=Rj
';RRRRRRRR1_mq)R t:HRL0=R:R''j;R
RRRRRRzRvppaqzXdn4vU_mR7 :MRH0CCos=R:R-j;-dj:nUG4R-+/RRB;4B:qBR/j+nRdG;4URR.:d4nGURR+BQq1
RRRRRRRRqB_717_z:ARR0LHRR:=';j'-'-RjR':N;88R4R''#:RkSL
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2R;
R
RRSsbF0
R5SRSq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSA:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;SRSB:MRHR8#0_oDFHPO_CFO0sd56RI8FMR0Fj
2;S1SqQ,thRQA1tRh,qpBBmRq7:MRHR8#0_oDFH
O;S SBRH:RM0R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
S1BqQRR:H#MR0D8_FOoH_OPC05Fs68cRF0IMF2Rj;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;S
SBmq1RF:Rk#0R0D8_FOoH_OPC05Fs68cRF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpqdpznUX4RB:RFFlbM0CMRRH#0Csk;R
RR-R
-------------------------v--zqpa7p7qzX4U4-U--------------------------------------m
Bvhum Rhavazpqq77pUz4X
4USMoCCOsH5S
Sq j)tRR:LRH0:'=Rj-';-jR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
ASSjt) RL:RH:0R=jR''
;RS4Sq)R t:HRL0=R:R''j;S
SA 4)tRR:LRH0:'=Rj
';S)SB :tRR0LHRR:=';j'
mSSz)a_ :tRR0LHRR:=';j'
uSSQju _t) RL:RH:0R=jR''S;
SuuQ )4_ :tRR0LHRR:=';j'
qSS1hQtj _)tRR:LRH0:'=Rj
';S1SAQjth_t) RL:RH:0R=jR''S;
SQq1t_h4)R t:HRL0=R:R''j;S
SAt1Qh)4_ :tRR0LHRR:=';j'
qSSBmBpq)7_ Rtj:HRL0=R:R''j;S
SqpBBm_q7)4 tRL:RH:0R=jR''R;
RRRRR1RRm)q_ :tRR0LHRR:=';j'
ASS_7q7_A1zRL:RH:0R=jR''R;R-'-RjR':N;88R''4:kR#LS
SB7_q7z_1ARR:LRH0:'=Rj
';SzSvp7aq7zqp44UXUm_v7: RR0HMCsoCRR:=j-;-jU:4GR4U+R/-44UGU/R+-;RBR:R4RBqB/+jRRG4U4+UR/4-RUUG4;:R.44UGU/R+-UR4GR4U+qRB1SQ
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5SjSq,Rq4:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SjSA,RA4:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SQS1qQ,1ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S
SBRR:H#MR0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R
RRRRRR1RqQ,thAt1QhRR:H#MR0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RRRRRRRR q1p1,A :pRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;R
RRRRRRqRB1:QRRRHM#_08DHFoOC_POs0F5R6c8MFI0jFR2R;
RRRRRqRRBmBpq:7RRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R
RRRRRRmR1qm,1ARR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
S1BqmRR:FRk0#_08DHFoOC_POs0F5R6c8MFI0jFR22
S;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvza7q7q4pzUUX4RB:RFFlbM0CMRRH#0Csk;-

-------------------------v--zqpapUz4X-4U-------------------------------------B-
mmvuha hRpvzazqp44UXUo
SCsMCH
O5S)Sq :tRR0LHRR:=';j'-'-RjR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCS
SAt) RL:RH:0R=jR''
;RS)SB :tRR0LHRR:=';j'
7SS)R t:HRL0=R:R''j;R
RRRRRRzRma _)tRR:LRH0:'=Rj
';SQSuu) _ :tRR0LHRR:=';j'
qSS1hQt_t) RL:RH:0R=jR''S;
SQA1t)h_ :tRR0LHRR:=';j'
7SS1hQt_t) RL:RH:0R=jR''S;
SBqBp7mq_t) jRR:LRH0:'=Rj
';SBSqBqpm7 _)t:4RR0LHRR:=';j'
ASS_7q7_A1zRL:RH:0R=jR''R;R-'-RjR':N;88R''4:kR#LS
SB7_q7z_1ARR:LRH0:'=Rj
';SzSvppaqzX4U4vU_mR7 :MRH0CCos=R:R-j;-qj:BjB/R-+/RG4U4+UR/B-R;:R4q/BBj/R+-UR4GR4U+qRB1RQ;.4:RUUG4R-+/R+7RR1BqQS;
Spvza _)1_ av m7R#:R0MsHo=R:RY"1hRB"-1-RY,hBRYq1hSB
2
;
SsbF0
R5SRSq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;SRSA:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;S,SBR:7RRRHM#_08DHFoOC_POs0F5R6d8MFI0jFR2R;
RRRRRqRR1hQt,1RAQRth:MRHR8#0_oDFH
O;RRRRRRRRBQq1RH:RM0R#8F_Do_HOP0COF6s5cFR8IFM0R;j2
RRRRRRRRBqBp7mq,Q71t:hRRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;S
SBmq1RF:Rk#0R0D8_FOoH_OPC05Fs68cRF0IMF2Rj
;S2
7 hRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVvazpq4pzUUX4RB:RFFlbM0CMRRH#0Csk;-

-------------------------q--pcz67------------------------------------
--Bumvmhh apRqz76c
CSoMHCsOS5
RRRRqt) RL:RH:0R=jR''-;R-''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8CRRRRRRRRAt) RL:RH:0R=jR''S;
RRRRqt1Qh _)tRR:LRH0:'=Rj
';SRRRRQA1t)h_ :tRR0LHRR:=';j'
RSRRBRqBqpm7 _)tRR:LRH0:'=Rj
';SRRRRamz_t) RL:RH:0R=jR''S;
RRRRA7_q7z_1ARR:LRH0:'=Rj-';-''j:8N8;4R''k:#LR
SRBRR_7q7_A1zRL:RH:0R=jR''R;
RRRRRqRRp_z7v m7RH:RMo0CC:sR=;Rj-:-jq/BBj/R+-RRA+R/-q4;R:BqB/+jR/A-RRB+Rq;1QRq.:R-+/R+ARR1BqQS;
Szqp_1)  va_mR7 :0R#soHMRR:="h1YB-"R-h1YBq,R1BYh
RRRR
2;RRRRb0FsRS5
RRRRqRR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRARR:H#MR0D8_FOoH_OPC0RFs5R6d8MFI0jFR2S;
RRRRB: RRRHM#_08DHFoOS;
RRRRBRpi:MRHR8#0_oDFH
O;SRRRR1)  :aRRRHM#_08DHFoOS;
RRRRqt1Qh1,AQRth:MRHR8#0_oDFH
O;SRRRRBqBp7mqRH:RM0R#8F_Do;HO
RSRRqRB1:QRRRHM#_08DHFoOC_POs0FRc56RI8FMR0Fj
2;SRRRRz7maRR:FRk0#_08DHFoOC_POs0FRd56RI8FMR0Fj
2;SRRRR1BqmRR:FRk0#_08DHFoOC_POs0FRc56RI8FMR0FjR2
R2RR;h
 7mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzqp6Rc7:FRBlMbFCRM0H0#Rs;kC
-
------------------------------p-up------------------------
--Bumvmhh apRupR
RR RthQ )BR5
RRRRRRRRRRRRwiBpQ:hRR)1aQRht:"=R43jjjR";-s-VCCJkMRO$F0VREOCRDM	H5
v2RRRRRRRRRRRRRe7 QRB :aR1)tQhRR:=".tWqU-4"-;R-W"t.4q-U"",tqW.-"66,W"t.-q)4
U"RRRRRRRRRRRRRh7Y_QQ7e _1pRR:1Qa)h:tR=VR"NCD#"-;-0Csk:1Q7 Rp;V#NDC7:QQ1e_ Rp
RRRRRRRRRRRRQe7Q_p1 RH:RMo0CC:sR=;Rj-M-QbRk08HHP8RCsQe7Q,:Rj4:,4.333nnd:cR3R4c~n
RRRRRRRRRRRRYR7hA_w7_Qe1R p:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRARw7_Qe1R p:MRH0CCos=R:R-j;-CwC8OLN	HR8PCH8sARw7,QeR:Rj4:,4.333nnd:c43R~
ncRRRRRRRRRRRRRh7Y_Qm7e _1pRR:1Qa)h:tR=VR"NCD#"-;-0Csk:1m7 Rp;V#NDC7:mQ1e_ Rp
RRRRRRRRRRRRme7Q_p1 RH:RMo0CC:sR=;RU-/-.c//U4dn/.U/c//ncUgj/n4/4../4UR
RRRRRRRRRRuRR1_7q1R p:aR1)tQhRR:="jjjj-";-R
RRRRRRRRRR7RRY7h_qh_ R1:Rah)Qt=R:RN"VD"#C;0--s:kCuq17RRFs7Yza7FqRs7RwqV;RNCD#:qR7_p1 
RRRRRRRRRRRRzR7aqY7_p1 R1:Rah)Qt=R:Rj"4j;j"-R-
RRRRRRRRRRRRBmpizwa_aQ_7)RR:LRH0:'=R4R';-B-RpzimaHRVM0CRkMMHoHR8s0COH3FMR''4RDFM$R
RRRRRRRRRRBRRpzimawu_aQ_7)RR:LRH0:'=R4R';-'-R4F'RM
D$RRRRRRRRRRRRRiBpm_za7_pY1ua RH:RMo0CC:sR=;RjRR--j,,4.
,cRRRRRRRRRRRRRiBpmuza_Y7p_ 1auRR:HCM0oRCs:j=R;-R-R4j,,
.
RRRRRRRRRRRRRiBpm7zad)_1BRR:1Qa)h:tR=BR"pzima-";-D#CCRO08dHPR0Fkb,k0RiBpmuzaRRFsBmpizRa
RRRRRRRRRRRRBwpiA _1pRR:1Qa)h:tR=HR"Ms0CM"ND;"--HCM0sDMN"C,"Gs0CM"ND
RRRRRRRRRRRRpRBiamz_uAYqR11:aR1)tQhRR:="DVN#;C"
RRRRRRRRRRRRpRBiamzuY_Au1q1R1:Rah)Qt=R:RN"VD"#C;R
RRRRRRRRRRBRRpzimaA7_Y1uq1RR:1Qa)h:tR=VR"NCD#"R;
RRRRRRRRRRRRBmpiz_a71R)B:aR1)tQhRR:="iBpm"za;#--CODC0HR8PkRF00bk,BRRpzimaFuRspRBiamz
RRRRRRRRRRRRYR7h7_1Q1e_ :pRR0HMCsoCRR:=.-R-R4.~.FU,MRD$CMPCRlMk
RRRRRRRRRRRRRR
RRRSRRRRR;R2
RRRR)umaR5
RRRRRRRRRRRRBQpihRR:Q#hR0D8_FOoH;R
RRRRRRRRRRBRRpAiwRQ:Rh0R#8F_Do:HO=''j;R
RRRRRRRRRRQRR7p1 RQ:RM0R#8F_Do_HOP0COF6s5RI8FMR0Fj
2;RRRRRRRRRRRRR7wA1R p:MRQR8#0_oDFHPO_CFO0sR568MFI0jFR2R;
RRRRRRRRRRRRm 71pRR:Q#MR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
RRRRRRRRRRRR R)1R a:MRHR8#0_oDFH=O:';j'
RRRRRRRRRRRR R)1_ auRR:H#MR0D8_FOoH:j=''R;
RRRRRRRRRRRR)  1aR_Q:RHM#_08DHFoO':=j
';RRRRRRRRRRRRR1)  1a_RH:RM0R#8F_DoRHO:j=''R;
RRRRRRRRRRRRuq17,pw7YRR:Q#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
RRRRRRRRRRRRzR7aqY7RQ:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;RRRRRRRRRRRRRBpmiRR:mRza#_08DHFoOR;
RRRRRRRRRRRRBmpiz:aRRamzR8#0_oDFH
O;RRRRRRRRRRRRRiBpm7zaRF:Rk#0R0D8_FOoH;R
RRRRRRRRRRBRRpzima:uRR0FkR8#0_oDFH
O;RRRRRRRRRRRRRiBpm7zadRR:FRk0#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVuRpp:FRBlMbFCRM0H0#Rs;kC
-
------------------------------p-Bie7Q-------------------------B-
mmvuha hRiBp7
QeRRRRt  h)5QB
RSRR7RRQve_mR7 :aR1)tQhRR:=";."RR--",."R3"d6R",",c"R""6
RSRRtRR1h) R1:Rah)Qt=R:RN"VD"#CRR--"DVN#,C"Rs"0k
C"SRRRR
2;RRRRuam)5R
RRRRRR]RRBQpihRR:Q#hR0D8_FOoH;R
SRRRR)  1a:hRRRQh#_08DHFoOS;
RRRRRpBqQ:ARRRQM#_08DHFoOS;
RRRRRiBpmRza:zRma0R#8F_Do
HORRRRRRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRBie7QRB:RFFlbM0CMRRH#0Csk;-

-----------------------------7--]hB -------------------------------------m
Bvhum Rha7 ]BhR
RRmRu)5aR
BSRpzimaRR:mRza#_08DHFoO
;SS RBRQ:Rh0R#8F_Do;HOSR
SBQpihRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7 ]BhRR:BbFlFMMC0#RHRk0sCR;RR

S-----------------17T---------------------------------m
Bvhum Rha7
T1RRRRt  h)5QB
RSRRQRwwvm_m_7 1R p:HRL0=R:R''j;R--wmQwR8lFCCR#D0CO:jR''7,7)CRll$FsR8lFC4;''t:R7R7)lCF8
)SS7h_ua:)RR0LH_OPC0RFs:"=Rj"jj;w--QRwms8CNRHbFMs0CR0#C0oHM
7SSTv1_mR7 :0R#soHMRR:=""X4;-R-R4"X"X,".7_7),.""_X.7d7)"X,"c"",X7._7_)d "Xa
RRRRRRRRp]WR#:R0MsHo=R:RN"VD"#C;"--0Csk"";RV#NDCR"
RSRRt 1)hRR:#H0sM:oR=VR"NCD#"-R-V#NDC0,Rs
kCS
2;RRRRuam)5R
RRRRRRTR71,QhuiBp,pwBi ,)1R a:MRHR8#0_oDFH
O;S S)q:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S)iBp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
Sp7p1ua ,aW1 :uRRRHM#_08DHFoOC_POs0F58(RF0IMF2Rj;S
S)qpm7Rh,)evm ),R7,Q)Rp]m7RR:H#MR0D8_FOoH;R
RRRRRRpRWmhq7,vRWm,e RQW7)RR:H#MR0D8_FOoH;R
RRRRRRTR71j)g,TR71,WjR17TWj.(RF:Rk#0R0D8_FOoH;S
S)QumhRa,WQumh:aRR0FkR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
Sq)ep,Q7))Az1Ra,)qwptW,RwtpqRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRT:1RRlBFbCFMMH0R#sR0k
C;
----------------------------7--ppp7Y---------------------------------------
vBmu mhh7aRppp7YR
RR RthQ )BR5
RRRRR7RRpQp_hp1 RL:RH:0R=jR''-;R-''j:bL$NR##lCF8,4R''k:R#8CRD8D_C$DNRDOCDR
RRRRRRpR7YQ_1t:hRR0LHRR:=';j'RR--':j'',+'R4R''':R-R'
RRRRR7RRpqY_7:KRR0HMCsoCRR:=j-R-j6~.68,RD#$_H=oMj8R:DN$_8R[;8_D$#MHo=R4:-n.6+$8D_[N8RR
RR;R2
RRRR)umaR5
RRRRR7RRpap1 :uRRRQh#_08DHFoOC_POs0F58(RF0IMF2Rj;R
RRRRRRpRBi:QhQ#hR0D8_FOoH;R
RRRRRRQR7)m,pq,7hv me:MRQR8#0_oDFH
O;RRRRRRRRBmpiz:aRRamzR8#0_oDFH
O;RRRRRRRRwtpqRm:Rz#aR0D8_FOoH
RRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV77ppp:YRRlBFbCFMMH0R#sR0k
C;RRRR
--------------------------------17B-------------------------------------m
Bvhum Rha7
B1RRRRt  h)RQB5S
S7_B1v m7R#:R0MsHo=R:RQ")1tQh"RRR-p-BiBj,p,i4B.pi,iBpdh,t7B,eBQ,)1tQh,pwqptQh,iBpjh_t7p,Biej_BBB,p_i4t,h7B4pi_BeB,iBp.h_t7p,Bie._BBB,p_idt,h7Bdpi_BeB
;S2
mSu)5aR
BSSpRij:hRQR8#0_oDFH
O;SpSBi:4RRRQh#_08DHFoOS;
SiBp.RR:Q#hR0D8_FOoH;S
SBdpiRQ:Rh0R#8F_Do;HO
BSSp i1pRR:Q#hR0D8_FOoH_OPC05FsdFR8IFM0R;j2
1SS mpw)RB :hRQR8#0_oDFH
O;SpSBiamzRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7RB1:FRBlMbFCRM0H0#Rs;kCRRRR
-
------------------------------T-7B- ----------------------------------
--Bumvmhh aTR7BR 
RuRRmR)a5R
SBmpiz:aRRamzR8#0_oDFHSO;
BSR RR:Q#hR0D8_FOoH;SS
RiBpQ:hRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRB7T RR:BbFlFMMC0#RHRk0sCR;RRRR
RCR
MO8RFFlbM0CM#R;RR
R

