--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb/oIlbNbC/s#GHHDMDG/HoL/CsMCHoO/CoM_CsMCHsO/Nsl_IE3P8Ry4f-
-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00X$R)4qv.4UX1#RH
bRRFRs05R
RRRRRRRRmRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.RRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcRRR:H#MR0k8_DHFoOR;
RRRRRqRR6RRR:MRHR8#0_FkDo;HO
qSSnRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RRH:RM0R#8D_kFOoH;R
RRRRRRBRWp:iRRRHM#_08koDFH
O;RRRRRRRRWR RRH:RM0R#8D_kFOoH
RRRRRRR2C;
MX8R)4qv.4UX1
;
NEsOHO0C0CksRv)q_FeRV)RXq.v4U1X4R
H##MHoN0DRj0,R4RR:#_08koDFH
O;#MHoNIDRCR4,IRC.:0R#8D_kFOoH;C
Lo
HMRRRRRRRRRRRRXqz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,6RqRR=>q
6,SSSSSRSRW= R>CRI4W,RBRpi=W>RB,piR=mR>jR02R;
RRRRRRRRRXRR4qz)vRnc:qR)vXnc4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,6RqRR=>q
6,SSSSSRSRW= R>CRI.W,RBRpi=W>RB,piR=mR>4R02m;
RR<=0IjRERCMq=nRR''jR#CDC4R0;C
I4=R<RRW NRM8M5F0q;n2
.ICRR<=WN RMq8Rn
;
CRM8)_qve
;

LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$)RXqcvnXR.1HR#
RsbF0
R5RRRRRRRRmRjRRF:Rk#0R0k8_DHFoOR;
RRRRRmRR4RRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4RRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq6RRR:H#MR0k8_DHFoOR;
RRRRR7RRjRRR:MRHR8#0_FkDo;HO
RRRRRRRRR74RRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpi:MRHR8#0_FkDo;HO
RRRRRRRRRW RRR:H#MR0k8_DHFoOR
RRRRRR
2;CRM8Xv)qn.cX1
;
NEsOHO0C0CksRv)qn.cX1R_eFXVR)nqvc1X.R
H#LHCoMR
RRRRRRRRRRzRX)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R,7jRRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qcRRq6=q>R6S,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,RRR=>m;j2
RRRRRRRRRRRRzX4)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R,74RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qcRRq6=q>R6S,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,RRR=>m;42
8CMRv)qn.cX1;_e
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00X$R)dqv.1XUR
H#RFRbs50R
mSSRF:Rk#0R0D8_FOoH_OPC05FsR8(RF0IMF2Rj;R
RRRRRRjRqR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRH:RM0R#8D_kFOoH;R
RRRRRR.RqR:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRH:RM0R#8D_kFOoH;R
RRRRRRcRqR:RRRRHM#_08koDFH
O;RRRRRRRR7RRRRH:RM0R#8F_Do_HOP0COF5sRR8(RF0IMF2Rj;R
RRRRRRBRWp:iRRRHM#_08koDFH
O;RRRRRRRRWR RRH:RM0R#8D_kFOoH
RRRRRRR2C;
MX8R)dqv.1XU;N

sHOE00COkRsC)_qveVRFRqX)vXd.UH1R#C
Lo
HMRRRRRRRRRRRRXqz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>5R7jR2,7>4=R4752q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rc
,RSSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m=jR>5RmjR2,m=4R>5Rm4;22
RRRRRRRRRRRRzX4)Rqv:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>725.,4R7=7>R5,d2RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qc
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRRmj=m>R5,.2RRm4=m>R52d2;R
RRRRRRRRRR.RXzv)qR):Rq.vdXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=Rc7527,R4R=>7256,jRqRR=>qRj,q=4R>4Rq,.RqRR=>q
.,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>qRd,q=cR>cRq,S
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,jRmRR=>m25c,4RmRR=>m2562R;
RRRRRRRRRXRRdqz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>5R7nR2,7>4=R(752q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>RcS,
SSSSSWRR >R=R,W RpWBi>R=RpWBim,Rj>R=Rnm52m,R4>R=R(m52
2;CRM8)_qveD;
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
M
C0$H0RqX)vXd.cH1R#R
Rb0FsRR5
RSRRm:jRR0FkR8#0_FkDo;HO
RRRR4SmRF:Rk#0R0k8_DHFoOR;
RSRRm:.RR0FkR8#0_FkDo;HO
RRRRdSmRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRH:RM0R#8D_kFOoH;R
RRRRRR4RqR:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRH:RM0R#8D_kFOoH;R
RRRRRRdRqR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRH:RM0R#8D_kFOoH;R
RR7RSjRRR:MRHR8#0_FkDo;HO
RRRR4S7R:RRRRHM#_08koDFH
O;RRRRSR7.RRR:H#MR0k8_DHFoOR;
RSRR7RdRRH:RM0R#8D_kFOoH;R
RRRRRRBRWp:iRRRHM#_08koDFH
O;RRRRRRRRWR RRH:RM0R#8D_kFOoH
RRRRRRR2C;
MX8R)dqv.1Xc;N

sHOE00COkRsC)_qveVRFRqX)vXd.cH1R#C
Lo
HMRRRRRRRRRRRRXqz)vRR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>jR7,4R7=7>R4q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=R,qdRRqc=q>Rc
,RSSSSSRSRW= R> RW,BRWp=iR>BRWpRi,m=jR>jRm,4RmRR=>m;42
RRRRRRRRRRRRzX4)Rqv:qR)vXd..
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>7R.,7>4=R,7dRRqj=q>Rjq,R4>R=R,q4RRq.=q>R.R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=q>Rdq,Rc>R=R,qc
SSSSRSSRRW =W>R W,RBRpi=W>RB,piRRmj=m>R.m,R4>R=R2md;M
C8qR)v;_e
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3ND
;
CHM00X$R)4qvn1XUR
H#RFRbs50R
mSSRF:Rk#0R0D8_FOoH_OPC0RFs5RR(8MFI0jFR2R;
RRRRRqRRjRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4RRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRR:MRHR8#0_oDFHPO_CFO0sRR5(FR8IFM0R;j2
RRRRRRRRpWBiRR:H#MR0k8_DHFoOR;
RRRRRWRR RRR:MRHR8#0_FkDo
HORRRRR2RR;M
C8)RXqnv4X;U1
s
NO0EHCkO0s)CRqev_RRFVXv)q4UnX1#RH
oLCHRM
RRRRRRRRRXRRzv)qR):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5j>R=Rj7527,R4R=>7254,.R7RR=>725.,dR7RR=>725d,SR
SRSSRRRRRRRRRRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qdRS
SSSSSR RWRR=>WR ,WiBpRR=>WiBp,SR
SSSSSmRRj>R=Rjm52m,R4>R=R4m52m,R.>R=R.m52m,Rd>R=Rdm52
2;RRRRRRRRRRRRX)4zq:vRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=7>R5,c2R=74>5R76R2,7=.R>5R7nR2,7=dR>5R7(R2,
SSSSRRRRRRRRqRRj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>Rd
,RSSSSSRSRW= R> RW,BRWp=iR>BRWpRi,
SSSSRSSRRmj=m>R5,c2RRm4=m>R5,62RRm.=m>R5,n2RRmd=m>R52(2;M
C8qR)v;_e

-----
-HR1lCbDRv)qR0IHEHR#MCoDR7q7)1 1RsVFR0LFECRsNN8RMI8RsCH0
R--aoNsC:0RRDXHH
MG-D-
HNLssH$RC;CC
Ck#RCHCC03#8F_Do_HO4c4n3DND;#
kCCRHC#C30D8_FOoH_o#HM3C8N;DD
LDHs$NsRHkM#;Hl
Ck#RHkM#3HlPlOFbCFMM30#N;DD
0CMHR0$)_qv)HWR#R
RRCRoMHCsO
R5RRRRRRRRVHNlD:$RRs#0HRMo:"=RMCFM"R;
RRRRRIRRHE80RH:RMo0CC:sR=;RURR
RRRRRR8RN8HsI8R0E:MRH0CCos=R:RRU;RRRRR-RR-HRLoMRCFEkoRsVFRb8C0RE
RRRRR8RRCEb0RH:RMo0CC:sR=6R.nR;
RRRRR8RRF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRR-E-RNF#Rkk0b0CRsoR
RRRRRRHR8MC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#NR80HNRM0bkRosC
RRRRRRRR8N8sC_soRR:LDFFCRNM:V=RNCD#RRRRR-R-R8ENR8N8s#C#RosC
RRRRRRRR
2;RRRRb0FsRR5
RRRRR7RRm:zaR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
RRRRRRRRh7QRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;
RRRRRqRR7R7):MRHR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRW RH:RM0R#8F_Do;HORRRRR-RR-sRIHR0CCLMNDVCRFssRNRl
RRRRRBRRp:iRRRHM#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
RRRRRRRRpmBiRR:H#MR0D8_FOoHRRRRR-RR-bRF0DROFRO	VRFs80Fk
RRRRRRRR
2;CRM8CHM00)$Rq)v_W
;
---
-HRwsR#0HDlbCMlC0HN0FlMRkR#0LOCRNCDD8sRNO
Ej-N-
sHOE00COkRsCLODF	N_slVRFRv)q_R)WH
#
ObFlFMMC0)RXq.v4U1X4
FRbs50R
RRRmRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRRq:6RRRHM#_08DHFoOR;
RnRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;


ObFlFMMC0)RXqcvnX
.1RsbF0
R5RmRRjRR:FRk0#_08DHFoOR;
R4RmRF:Rk#0R0D8_FOoH;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;RqRR6RR:H#MR0D8_FOoH;R
RRR7j:MRHR8#0_oDFH
O;R7RR4RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;O

FFlbM0CMRqX)vXd.cR1
b0FsRR5
RjRmRF:Rk#0R0D8_FOoH;R
RRRm4:kRF00R#8F_Do;HO
RRRm:.RR0FkR8#0_oDFH
O;RmRRdRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7:jRRRHM#_08DHFoOR;
R4R7RH:RM0R#8F_Do;HO
RRR7:.RRRHM#_08DHFoOR;
RdR7RH:RM0R#8F_Do;HO
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMMX0R)dqv.1XU
b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
F
OlMbFCRM0Xv)q4UnX1b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
VOkM0MHFRMVkOM_HHL05RL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
RRHV5RL20MEC
RRRR0sCk5sM";"2
CRRD
#CRRRRskC0s"M5BDFk8FRM0lRHblDCCRM0AODF	qR)vQ3R#ER0CCRsNN8R8C8s#s#RC#oH0CCs8#RkHRMo0REC#CNlRFODON	R#ER0CqR)v2?";R
RCRM8H
V;CRM8VOkM_HHM0V;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHoN;
0H0sLCk0RMoCC0sNFss_CsbF0VRFRFLDOs	_N:lRRONsECH0Os0kC#RHRMVkOM_HHN058_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+4-;
-MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R55580CbERR-4/2RR2d.R5+R5C58bR0E-2R4R8lFR2d.R4/Rn;22R-RR-RRyF)VRq.vdXR41ODCD#CRMC88CR-
-O#FM00NMRVDC0P_FC:sRR0HMCsoCRR:=5855CEb0R4+R6l2RFd8R./2RR24n;RRRRRRRRRRRRRRRRRRRRRRRR-R-RFyRVqR)vX4n4M1RCCC88FRVsCRDVF0RPRCsI8Fs#$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDF_k0s4CoR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFEROFCF#R0LCIMCCRh7QR8NMR0FkbRk0FAVRD	FORv)q
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7R7)VRFsI0sHCH
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoN)DRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7)q7#)
HNoMDqRW7_7)0Rlb:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMCW7q7)H
#oDMNRh7Q_b0lR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFHRbbHCDM7CRQ#h
HNoMD RW_b0lR#:R0D8_FOoH;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR
W -C-RML8RD	FORlsNRbHlDCClM00NHRFM#MHoN
D#
R--LHCoMCR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bRVDC0CFPsR_0HN#Rs$sNRR5j0dFR2VRFR0HMCsoC;$
0bDCRCFV0P_Cs0R_.HN#Rs$sNRR5j04FR2VRFR0HMCsoC;k
VMHO0FbMRNH85R#:R0D8_FOoH_OPC0;FsR,I4RRI.:MRH0CCoss2RCs0kM0R#8F_Do_HOP0COFHsR#N
PsLHNDPCRN:sRR8#0_oDFHPO_CFO0s45I-84RF0IMF2Rj;C
Lo
HMRFRVsRR[HPMRNss'NCMoRFDFbR
RRVRHRR5[<I=R.02RERCM
RSRP5Ns[:2R=5RHHF'DI2+[;C
SD
#CSPRRN[s52=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsMP;Ns
8CMR8bN;k
VMHO0FoMRCI0_HE80_IU5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0UE/;R
RH5VR58IH0lERFU8R2RR>c02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_U
MVkOF0HMCRo0H_I8_0E.H5I8:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=I0H8E;/.
sRRCs0kMNRPDC;
Mo8RCI0_HE80_
.;VOkM0MHFR0oC_8IH0IE5HE80RH:RMo0CCRs2skC0sDMRCFV0P_Cs0R_.HP#
NNsHLRDCPRND:CRDVP0FC0s__
.;LHCoMR
RP5ND4:2R=CRo0H_I8_0E.H5I820E;R
RH5VRI0H8EFRl8RR.=2RjRC0EMR
RRNRPD25jRR:=jR;
R#CDCR
RRNRPD25jRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCI0_HE80;k
VMHO0FoMRCI0_HE8058IH0:ERR0HMCsoC2CRs0MksRVDC0CFPsR_0HP#
NNsHLRDCPRND:CRDVP0FC0s_RR:=5Rj,jj,R,2Rj;C
Lo
HMRNRPD25dRR:=o_C0I0H8E5_UI0H8E
2;RNRO#5CRI0H8EFRl82RUR
H#RERICcMRRd|RRR=>P5ND.:2R=;R4
IRRERCM.>R=RDPN5R42:4=R;R
RIMECR=4R>NRPD25jRR:=4R;
RCIEM0RFE#CsRR=>MDkD;R
RCRM8OCN#;R
RskC0sPMRN
D;CRM8o_C0I0H8EO;
F0M#NRM0#H_I8_0ENNss$RR:D0CVFsPC_:0R=CRo0H_I850EI0H8E
2;O#FM00NMRI#_HE80_sNsNn$_cRR:D0CVFsPC_.0_RR:=o_C0I0H8EH5I820E;k
VMHO0FoMRCM0_k4l_.8U5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C04E/.
U;RVRHR855CEb0R8lFRU4.2RR>424.RC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._4UV;
k0MOHRFMo_C0D0CVFsPC_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF842.U;M
C8CRo0C_DVP0FCns_cV;
k0MOHRFMo_C0M_kln8c5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
RRRH5VR80CbE=R<R.44R8NMRb8C0>ERR2cURC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FC8s5CEb0RH:RMo0CCRs;lRNG:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E-NRlG=R>RRj20MEC
RRRRDPNRR:=80CbERR-l;NG
CRRD
#CRRRRPRND:8=RCEb0;R
RCRM8H
V;RCRs0Mks5DPN2C;
Mo8RCD0_CFV0P;Cs
MVkOF0HMCRo0k_Ml._d5b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=URcR8NMRb8C0>ERR24nRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;d.
MVkOF0HMCRo0k_Mln_45b8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0<ER=nR4R8NMRb8C0>ERRRj20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kl4
n;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88OR
F0M#NRM0M_klODCD_U4.RH:RMo0CC:sR=CRo0k_Ml._4UC58b20E;F
OMN#0MD0RCFV0P_Csn:cRR0HMCsoCRR:=o_C0D0CVFsPC_5nc80CbE
2;O#FM00NMRlMk_DOCDc_nRH:RMo0CC:sR=CRo0k_Mlc_n5VDC0CFPsc_n2O;
F0M#NRM0D0CVFsPC_Rd.:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCns_cn,Rc
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$C._4U#RHRsNsN5$RM_klODCD_U4.RI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_RncHN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._dRRH#NNss$MR5kOl_C_DDd8.RF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0b4C_n#RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk_U4.RF:RkL0_k0#_$_bC4;.URRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rnc:kRF0k_L#$_0bnC_cR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kd#_.RR:F_k0L_k#0C$b_;d.RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_R4n:kRF0k_L#$_0b4C_nR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoN#DR_0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DD4R.U8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CnM_cRR:#_08DHFoO#;
HNoMDkRF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDF_k0C4M_nRR:#_08DHFoO#;
HNoMD_R#I_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_OD4D_.8URF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CnM_cRR:#_08DHFoO#;
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMD_R#HsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoN#DR_0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRND#8_N_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F58nRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2F
OMN#0MD0R#IL_HE80RH:RMo0CC:sR=HRI8-0EU#*5_8IH0NE_s$sN5-d24c2-*I#_HE80_sNsN.$52*-.#H_I8_0ENNss$254-I#_HE80_sNsNj$520;
$RbC0_lbNNss$HUR#sRNsRN$5I#_HE80_sNsNd$52R-48MFI0jFR2VRFR8#0_oDFHPO_CFO0sR5(8MFI0jFR2#;
HNoMDlR0b__UdR.,0_lbUn_4R0:RlNb_s$sNU-;
-MRC8CR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH

RRRcRzdRR:H5VRNs88_osC2CRoMNCs0-CR-CRoMNCs0LCRD	FORlsN
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRq&R757)j
2;RRRRRRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjj"jjRq&R757)4FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjj"jjRq&R757).FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjjjjjj&"RR7q7)R5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjj"jjRN&R8C_soR5d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjj&"RR7q7)R5c8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjRj"&8RN_osC58cRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRcR;
RzRR6:RRRRHV58N8s8IH0=ERRRn2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjj"jjRq&R757)6FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjj"jjRN&R8C_soR568MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjj"jjRq&R757)nFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjRj"&8RN_osC58nRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV58N8s8IH0=ERRRU2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jjjjj&"RR7q7)R5(8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjj&"RR7q7)R5U8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;R
RRMRC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjj"RR&q)7758gRF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=Rjjjj"RR&Ns8_Cgo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRNs88I0H8ERR=4R42oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"jRj"&7Rq74)5jFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&8RN_osC5R4j8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RRR:H5VRNs88I0H8ERR=4R.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR7q7)454RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<='Rj'&7Rq74)5.FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR''RR&Ns8_C4o5.FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=q)775R4d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=Ns8_C4o5dFR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
c;RRRRzR46RH:RVMR5F80RHsM_CRo2oCCMsCN0
RRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RCRRMo8RCsMCNR0Cz;46
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CR7)_mRzakM#Ho_R)miBp
RRRRnz4RRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soR42LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_so
4;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznR;
RzRR4R(R:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC4R;
RCRRMo8RCsMCNR0Cz;4(
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RsVFRHIs0kCR#oHMRiBp
RRRRUz4I:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0CzI4U;R
RR4Rzg:IRRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0Rgz4I
;
RRRR- -RGN0sRoDFHVORF7sRkRNDb0FsR#ONCR
RRsRzC:oRRFbsO#C#5iBp2CRLo
HMRRRRRVRHRp5Bie'  RhaNRM8BRpi=4R''02RE
CMRRRRR7RRQ0h_l<bR=QR7hR;
RRRRRqR)7_7)0Rlb<q=R7;7)
RRRRRRRW7q7)l_0b=R<R_N8s;Co
RRRRRRRW0 _l<bR= RW;R
RRRRRCRM8H
V;RRRRCRM8bOsFC;##
R
RR-R-RRQV)8CNR8q8s#C#RW=RsCH0R8q8s#C#,$RLb#N#Rh7QRR0FFbk0kH0RV RWRRH#CLMND
C8RRRRzGlkRb:RsCFO#W#5 l_0b),Rq)77_b0l,qRW7_7)0,lbRh7Q_b0l,kRF0C_soR2
RRRRRoLCHRM
RRRRRHRRVWR5q)77_b0lR)=Rq)77_b0lR8NMR_W 0Rlb=4R''02RE
CMRRRRRRRRRkRF0C_so<4R=QR7hl_0bR;
RRRRRCRRD
#CRRRRRRRRRkRF0C_so<4R=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRR8CMR;HV
RRRR8CMRFbsO#C#;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141R4
RzRR4:URRRHV5FOEH_OCI0H8ERR=4o2RCsMCN
0CRRRRRRRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
j;RRRR-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4z.;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRR.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vn_4dXUc4:7RRv)qA_4n114_4R
RRRRRRRRRRRRRRFRbsl0RN5bR75Qqj=2R>MRH_osC5,[2R7q7)=qR>FRDIN_I858s48dRF0IMF2Rj,QR7A>R=R""j,7Rq7R)A=D>RFsI_Ns885R4d8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25jRR=>F_k0L4k#5[H,2
2;
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
.;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1.1R.
RzRR.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CRRRRRRRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRR6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRd=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
6;RRRR-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRRnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rnz.;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRR.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..X7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_gU4.7X.R):Rq4vAn._1_
1.RRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co.+*[4FR8IFM0R[.*2q,R7q7)RR=>D_FII8N8s.54RI8FMR0FjR2,7RQA=">Rj,j"R7q7)=AR>FRDIN_s858s48.RF0IMF2Rj,R
RRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,RRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m5R42=F>RkL0_k5#.H*,.[2+4,mR7A25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC.Rz(R;
RRRRRCRRMo8RCsMCNR0Cz;.c
RRRR8CMRMoCC0sNC.RzdR;R
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cR
RR.RzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0RC
RRRRRzRR.:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNCdRzjR;
R-RR-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d4
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRRdRz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qvcnjgXRc7:qR)vnA4__1c1Rc
RRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7R)q=D>RFII_Ns885R448MFI0jFR27,RQ=AR>jR"j"jj,7Rq7R)A=D>RFsI_Ns885R448MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25dRR=>F_k0Lck#5RH,c+*[dR2,75mA.=2R>kRF0k_L#Hc5,[c*+,.2RR
RRRRRRRRRRRRRRmR7A254RR=>F_k0Lck#5cH,*4[+27,RmjA52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRRRRR8CMRMoCC0sNCdRz.R;
RRRRRCRRMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
RRRRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gRRRRzRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
RRRRRRRRczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRRdRz6RR:H5VRNs88I0H8ERR>4R42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d6
RRRRR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRRdRznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNCdRznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_.cUUX7RR:)Aqv41n_gg_1
RRRRRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7R)q=D>RFII_Ns885R4j8MFI0jFR27,RQ=AR>jR"jjjjj"jj,7Rq7R)A=D>RFsI_Ns885R4j8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm(A52>R=R0Fk_#LkU,5HU+*[(R2,75mAn=2R>kRF0k_L#HU5,[U*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A256RR=>F_k0LUk#5UH,*6[+27,RmcA52>R=R0Fk_#LkU,5HU+*[cR2,75mAd=2R>kRF0k_L#HU5,[U*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25.RR=>F_k0LUk#5UH,*.[+27,Rm4A52>R=R0Fk_#LkU,5HU+*[4R2,75mAj=2R>kRF0k_L#HU5,[U*2R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQ5uqj=2R>MRH_osC5[g*+,U2Ru7QA>R=R""j,mR7u=qR>bRFCRM,7Amu5Rj2=b>RN0sH$k_L#HU5,2R[2R;
RRRRRRRRRRRRRFRRks0_Cgo5*R[2<F=RkL0_k5#UH*,U[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[4<2R=kRF0k_L#HU5,[U*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R.2<F=RkL0_k5#UH*,U[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+dRR<=F_k0LUk#5UH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*c[+2=R<R0Fk_#LkU,5HU+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[6<2R=kRF0k_L#HU5,[U*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rn2<F=RkL0_k5#UH*,U[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+(RR<=F_k0LUk#5UH,*([+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*U[+2=R<RsbNH_0$LUk#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d(
RRRRRRRR8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
RRRRRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1_4U1
4URRRRzRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCR
RRRRRRdRzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRRc:jRRRHV58N8s8IH0>ERR24jRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRCRM8oCCMsCN0Rjzc;R
RR-R-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRRRRRzRRc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
4;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRRRRR.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qv4cj.X74nR):Rq4vAn4_1U4_1UR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7R)q=D>RFII_Ns8858gRF0IMF2Rj,QR7A>R=Rj"jjjjjjjjjjjjjj,j"R7q7)=AR>FRDIN_s858sgFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m5246RR=>F_k0L4k#n,5H4[n*+246,mR7Ac542>R=R0Fk_#Lk4Hn5,*4n[c+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rd2=F>RkL0_kn#454H,n+*[4,d2RA7m524.RR=>F_k0L4k#n,5H4[n*+24.,mR7A4542>R=R0Fk_#Lk4Hn5,*4n[4+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4Rj2=F>RkL0_kn#454H,n+*[4,j2RA7m5Rg2=F>RkL0_kn#454H,n+*[gR2,75mAU=2R>kRF0k_L#54nHn,4*U[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA(=2R>kRF0k_L#54nHn,4*([+27,RmnA52>R=R0Fk_#Lk4Hn5,*4n[2+n,mR7A256RR=>F_k0L4k#n,5H4[n*+,62RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A25cRR=>F_k0L4k#n,5H4[n*+,c2RA7m5Rd2=F>RkL0_kn#454H,n+*[dR2,75mA.=2R>kRF0k_L#54nHn,4*.[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4=2R>kRF0k_L#54nHn,4*4[+27,RmjA52>R=R0Fk_#Lk4Hn5,*4n[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Co4[U*+R4(8MFI04FRU+*[4,n2Ru7QA>R=Rj"j"R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmRuq=F>Rb,CMRu7mA254RR=>bHNs0L$_kn#45RH,.+*[4R2,7Amu5Rj2=b>RN0sH$k_L#54nH.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
.;RRRRRRRRCRM8oCCMsCN0Rgzd;R
RRMRC8CRoMNCs0zCRd
U;
RRRRRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dRn
RzRRdRUN:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNCR
RRRRRRdRzg:NRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRRRRRzRRcRjN:VRHR85N8HsI8R0E>2RgRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRc;jN
RRRRR--Q5VRNs88I0H8E=R<RRg2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4zcNR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRR)RAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7QRR=>"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR",q)77A>R=RIDF_8sN8Us5RI8FMR0Fj
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm=qR>bRFCRM,75mAdR42=F>RkL0_k.#d5dH,.+*[d,42RA7m52djRR=>F_k0Ldk#.,5Hd[.*+2dj,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5g=2R>kRF0k_L#5d.H.,d*.[+gR2,75mA.RU2=F>RkL0_k.#d5dH,.+*[.,U2RA7m52.(RR=>F_k0Ldk#.,5Hd[.*+2.(,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7An5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm.A56=2R>kRF0k_L#5d.H.,d*.[+6R2,75mA.Rc2=F>RkL0_k.#d5dH,.+*[.,c2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR7A.5.2>R=R0Fk_#LkdH.5,*d.[.+.27,Rm.A54=2R>kRF0k_L#5d.H.,d*.[+4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rj2=F>RkL0_k.#d5dH,.+*[.,j2RA7m524gRR=>F_k0Ldk#.,5Hd[.*+24g,mR7AU542>R=R0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5(=2R>kRF0k_L#5d.H.,d*4[+(R2,75mA4Rn2=F>RkL0_k.#d5dH,.+*[4,n2RA7m5246RR=>F_k0Ldk#.,5Hd[.*+246,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ac542>R=R0Fk_#LkdH.5,*d.[c+427,Rm4A5d=2R>kRF0k_L#5d.H.,d*4[+dR2,75mA4R.2=F>RkL0_k.#d5dH,.+*[4,.2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A4542>R=R0Fk_#LkdH.5,*d.[4+427,Rm4A5j=2R>kRF0k_L#5d.H.,d*4[+jR2,75mAg=2R>kRF0k_L#5d.H.,d*g[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mAU=2R>kRF0k_L#5d.H.,d*U[+27,Rm(A52>R=R0Fk_#LkdH.5,*d.[2+(,mR7A25nRR=>F_k0Ldk#.,5Hd[.*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7A256RR=>F_k0Ldk#.,5Hd[.*+,62RA7m5Rc2=F>RkL0_k.#d5dH,.+*[cR2,75mAd=2R>kRF0k_L#5d.H.,d*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>kRF0k_L#5d.H.,d*.[+27,Rm4A52>R=R0Fk_#LkdH.5,*d.[2+4,mR7A25jRR=>F_k0Ldk#.,5Hd[.*2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,7AQuRR=>"jjjjR",7qmuRR=>FMbC,mR7udA52>R=RsbNH_0$Ldk#.,5Hc+*[dR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA25.RR=>bHNs0L$_k.#d5cH,*.[+27,Rm5uA4=2R>NRbs$H0_#LkdH.5,[c*+,42Ru7mA25jRR=>bHNs0L$_k.#d5cH,*2[2;R
RRRRRRRRRRRRRRkRF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.zcNR;
RRRRRCRRMo8RCsMCNR0CzNdg;R
RRMRC8CRoMNCs0zCRd;UN
CRRMo8RCsMCNR0Cz;cd
zRRcRc:H5VRMRF0Ns88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<(#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jjjjj&"RRN#_8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj"jjR#&R__N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj&"RRN#_8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jRj"&_R#Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
cSzSH:RVNR58I8sHE80R6=R2CRoMNCs0SC
SIDF_8N8s=R<Rj"j"RR&#8_N_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;SSz6:VRHR85N8HsI8R0E=2RnRMoCC0sNCS
SD_FINs88RR<='Rj'&_R#Ns8_C6o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<#=R__N8s5ConFR8IFM0R;j2
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR(RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRRH#_MC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRR#M_H_osCRR<=7;Qh
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRzgRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=#k_F0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<#=R_0Fk_osC;R
RRMRC8CRoMNCs0zCR4
j;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz4:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRR#8_N_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz4R;
RzRR4:.RRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRR#8_N_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4
.;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4d:FRVsRRHH5MRM_klODCD_U4.R4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcz4RH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRR#RR_0Fk_5CMH<2R=4R''ERIC5MR#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRR_R#I_s0CHM52=R<RRW IMECR_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rcz4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4Rz6RR:H5VRNs88I0H8E=R<RR(2oCCMsCN0
RRRRRRRRRRRRRRRRF#_kC0_M25HRR<=';4'
RRRRRRRRRRRRRRRRI#_sC0_M25HRR<=W
 ;RRRRRRRRCRM8oCCMsCN0R6z4;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:nRRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qv.:URRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*.RU2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H442*.RU,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.v4URR:Xv)q4X.U4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5Co[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6R2,q=nR>FRDI8_N8ns52S,
SSSSSWRR >R=RI#_sC0_M25H,BRWp=iR>pRBim,RRR=>F_k0L_k#45.UH2,[2R;
RRRRRRRRRRRRR#RR_0Fk_osC5R[2<F=RkL0_k4#_.HU5,R[2IMECR_5#F_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRMRC8CRoMNCs0zCR4Rd;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR(z4RH:RVMR5kOl_C_DDn=cRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4RzU:NRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4NR;
RRRRRzRR4RUL:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_U4.Rj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECR#55__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UL
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRgz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4g
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_.:VRHR_5#I0H8Es_Ns_N$n4c52RR>jo2RCsMCN
0CRRRRRRRRzR.j:FRVsRR[H5MR#H_I8_0ENNss$c_n5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*-[RRR.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERR[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R54>R=RH#_MC_soH5I8-0E.-*[4R2,7=jR>_R#HsM_CIo5HE80-[.*-,.2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62
SSSSRSSRRW =I>RsC0_Mc_n,BRWp=iR>pRBim,R4>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4,jRmRR=>F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-2.2;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.[2-4RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-[.*-R.2<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[.I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNC.RzjS;
SMRC8CRoMNCs0zCRO_E	.S;
SORzE4	_RH:RV#R5_8IH0NE_s$sN_5ncj>2RRRj2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERR#.*_8IH0NE_s$sN_5nc4-2RRR42& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERR#.*_8IH0NE_s$sN_5nc4;22
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_soH5I8-0E._*#I0H8Es_Ns_N$n4c522-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,S
SSSSSR RWRR=>I_s0CnM_cW,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.#H_I8_0ENNss$c_n5-424;22
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#.*_8IH0NE_s$sN_5nc442-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.#H_I8_0ENNss$c_n5-424I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNCORzE4	_;R
SRRRRCRM8oCCMsCN0R(z4;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:4RRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN..RH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.N
RRRRRRRR.z.LRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_c=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.LR;
RRRRRzRR.R.O:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
O;RRRRRRRRz8..RH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDc_n2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDc_n2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
8;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.d:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RW;R
RRRRRRMRC8CRoMNCs0zCR.
d;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:URRRHV5I#_HE80_sNsNd$52RR>jo2RCsMCN
0CSOSzED	_C:6RRRHV58IH0>ER=*RU#H_I8_0ENNss$25dR8NMR8IH0>ER=2RURMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.jH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R[-R*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-[R5-*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_soH5I8-0ED_#LI0H8E*-U[R+(8MFI0IFRHE80-LD#_8IH0UE-*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=Rb0l_dU_.25[2S;
SRSRR#RN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.H,I8-0ED_#LI0H8E*-U[[+H2=R<Rb0l_dU_.25[52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbU._d5I#_HE80_sNsNd$522-42S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Ud#.5_8IH0NE_s$sN5-d24H25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d2.FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C5*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so*5U[R+(8MFI0UFR*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=Rb0l_dU_.25[2S;
SNSS#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdU.,*H[+[<2R=lR0b__Ud[.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CUo5*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloUC52R;
RRRRRRRRRRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_.25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d55j2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHR_5#I0H8Es_Ns5N$.>2RRRj2oCCMsCN0
RRRRRRRRcz._:cRRRHV58IH0>ER=2RcRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>_R#HsM_Cdo527,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,
SSSSRSSRRmd=F>RkL0_kd#_.k5MlC_ODdD_.2,d,.RmRR=>F_k0L_k#dM.5kOl_C_DDd..,2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.4R2,m=jR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Cod<2R=kRF0k_L#._d5lMk_DOCD._d,Rd2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_5d.M_klODCD_,d..I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_kd#_.k5MlC_ODdD_.2,jRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.cc_;R
RRRRRR.RzcR_d:VRHRH5I8R0E=2RdRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>jR''7,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_kd#_.k5MlC_ODdD_.2,.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDd4.,2m,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_5d.M_klODCD_,d..I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_kd#_.k5MlC_ODdD_.2,jRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.dc_;S
SCRM8oCCMsCN0REzO	;_c
zSSO_E	.RR:H5VR#H_I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRR.:cRRsVFRH[RM#R5_8IH0NE_s$sN5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>_R#HsM_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.R2,7=4R>_R#HsM_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[4R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
c;SMSC8CRoMNCs0zCRO_E	.S;
SEzO	R_4:VRHR_5#I0H8Es_Ns5N$j>2RRRj2oCCMsCN0
RRRRRRRRcz.RH:RVIR5HE80R8lFR=URRR42oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd.4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CojR2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,RRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
4;RRRRCRM8oCCMsCN0R4z.;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:6RRRHV5lMk_DOCDn_4R4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nN
RRRRRRRRnz.LRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.n;R
RRRRRR.Rzn:ORRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRNjRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.OR;
RRRRRzRR.Rn8:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
8;RRRRRRRRzC.nRH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RMR8R5N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzC.n;R
RRRRRR.Rzn:VRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.VR;
RRRRRzRR.Rno:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
o;RRRRRRRRzE.nRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
E;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.(:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRMRC8CRoMNCs0zCR.
(;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:URRRHV5I#_HE80_sNsNd$52RR>jo2RCsMCN
0CSOSzED	_C:6RRRHV58IH0>ER=*RU#H_I8_0ENNss$25dR8NMR8IH0>ER=2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Hn,[<2R=lR0b__U4jn52[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RM_R#I0H8Es_Ns5N$d42-RI8FMR0F4CRoMNCs0RC
RRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R[-R*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R5-R[2-4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)4qvnRR:Xv)q4UnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoI0H8E#-DLH_I8-0EU+*[HR[2<F=RkL0_k4#_nk5MlC_OD4D_nH,I8-0ED_#LI0H8E*-U[[+H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	C_D6S;
SEzO	0_o6RR:H5VRI0H8E=R>RNURMI8RHE80R8lFR>UR=2R6RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n_5#I0H8Es_Ns5N$d42-2
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54n#H_I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5U[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5[U*+8(RF0IMF*RU[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=Rb0l_4U_n25[2S;
SNSS#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Un,*H[+[<2R=lR0b__U4[n52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CUo5*H[+[<2R=kRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vR4n:)RXqnv4X
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbUn_452j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54njH25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;SMSC8CRoMNCs0zCRO_E	MS;
S8CMRMoCC0sNCORzEU	_;S
Sz	OE_:cRRRHV5I#_HE80_sNsN.$52RR>jo2RCsMCN
0CRRRRRRRRz_.gcRR:H5VRI0H8E=R>RRc2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>_R#HsM_Cdo527,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRS
SSSSSRdRmRR=>F_k0L_k#4Mn5kOl_C_DD4dn,2m,R.>R=R0Fk_#Lk_54nM_klODCD_,4n.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,,42RRmj=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rd2<F=RkL0_k4#_nk5MlC_OD4D_n2,dRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#n_45lMk_DOCDn_4,R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_54nM_klODCD_,4n4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.gcR;
RRRRRzRR.dg_RH:RVIR5HE80Rd=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>',j'RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>bRFCRM,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25.RR<=F_k0L_k#4Mn5kOl_C_DD4.n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R42<F=RkL0_k4#_nk5MlC_OD4D_n2,4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzg;_d
CSSMo8RCsMCNR0Cz	OE_
c;SOSzE.	_RH:RV#R5_8IH0NE_s$sN5R42>2RjRMoCC0sNCR
RRRRRRdRzjRR:VRFs[MRHR_5#I0H8Es_Ns5N$4-2RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-#U*_8IH0NE_s$sN5-d2.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4.nX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2RR74=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,42RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRRmj=F>RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R42<F=RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rjzd;S
SCRM8oCCMsCN0REzO	;_.
zSSO_E	4RR:H5VR#H_I8_0ENNss$25jRj>R2CRoMNCs0RC
RRRRRzRRd:4RRRHV58IH0lERFU8RR4=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CojR2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R4zd;S
SCRM8oCCMsCN0REzO	;_4
RRRRMRC8CRoMNCs0zCR.R6;RRRRRRRRRR
RR8CMRMoCC0sNCcRzcC;
MN8RsHOE00COkRsCLODF	N_sl
;
NEsOHO0C0CksR_MFsOI_E	CORRFV)_qv)HWR#F
OlMbFCRM0Xv)q4X.U4R1
b0FsRR5
RRRm:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
R6RqRH:RM0R#8F_Do;HO
RRRq:nRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
F
OlMbFCRM0Xv)qn.cX1b
RFRs05R
RRRmj:kRF00R#8F_Do;HO
RRRm:4RR0FkR8#0_oDFH
O;RqRRjRR:H#MR0D8_FOoH;R
RRRq4:MRHR8#0_oDFH
O;RqRR.RR:H#MR0D8_FOoH;R
RRRqd:MRHR8#0_oDFH
O;RqRRcRR:H#MR0D8_FOoH;R
RRRq6:MRHR8#0_oDFH
O;R7RRjRR:H#MR0D8_FOoH;R
RRR74:MRHR8#0_oDFH
O;RWRRBRpi:MRHR8#0_oDFH
O;RWRR RR:H#MR0D8_FOoH
;R2
8CMRlOFbCFMM
0;
lOFbCFMMX0R)dqv.1Xc
FRbs50R
RRRm:jRR0FkR8#0_oDFH
O;RmRR4RR:FRk0#_08DHFoOR;
R.RmRF:Rk#0R0D8_FOoH;R
RRRmd:kRF00R#8F_Do;HO
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RjR7RH:RM0R#8F_Do;HO
RRR7:4RRRHM#_08DHFoOR;
R.R7RH:RM0R#8F_Do;HO
RRR7:dRRRHM#_08DHFoOR;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0O;
FFlbM0CMRqX)vXd.U
1
RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRRq:cRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
ObFlFMMC0)RXqnv4X
U1RsbF0
R5RmRRRF:Rk#0R0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRq:jRRRHM#_08DHFoOR;
R4RqRH:RM0R#8F_Do;HO
RRRq:.RRRHM#_08DHFoOR;
RdRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
MVkOF0HMkRVMHO_M5H0LRR:LDFFC2NMR0sCkRsM#H0sMHoR#C
Lo
HMRVRHR25LRC0EMR
RRCRs0Mks5F"hRNsC8s/IHR0COVFMD0HORCOEOR	31kHlDHN0FlMRHN#l0ROEb#F#HCLDR"!!2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHRMVkOM_HHN058_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+4-;
-MOF#M0N0kRMlC_ODRD#:MRH0CCos=R:R55580CbERR-4/2RR2d.R5+R5C58bR0E-2R4R8lFR2d.R4/Rn;22R-RR-RRyF)VRq.vdXR41ODCD#CRMC88CR-
-O#FM00NMRVDC0P_FC:sRR0HMCsoCRR:=5855CEb0R4+R6l2RFd8R./2RR24n;RRRRRRRRRRRRRRRRRRRRRRRR-R-RFyRVqR)vX4n4M1RCCC88FRVsCRDVF0RPRCsI8Fs#$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lkd0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*RcI0H8Ek_MlC_OD+D#dFR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$Ldk#.RR:bHNs0L$_k.#d_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDF_k0s4CoR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFEROFCF#R0LCIMCCRh7QR8NMR0FkbRk0FAVRD	FORv)q
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7R7)VRFsI0sHCH
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8sN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRNDD_FII8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--I8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNsDRNs88_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2-;
-MRC8DRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD
#
-L-RCMoHRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMD0#
$RbCD0CVFsPC_H0R#sRNsRN$50jRF2RdRRFVHCM0o;Cs
b0$CCRDVP0FC0s__H.R#sRNsRN$50jRF2R4RRFVHCM0o;Cs
MVkOF0HMNRb8R5H:0R#8F_Do_HOP0COFRs;IR4,I:.RR0HMCsoC2CRs0MksR8#0_oDFHPO_CFO0s#RH
sPNHDNLCNRPsRR:#_08DHFoOC_POs0F5-I44FR8IFM0R;j2
oLCHRM
RsVFRH[RMNRPsN'sMRoCDbFF
RRRRRHV5<[R=.RI2ER0C
MRSPRRN[s52=R:RHH5'IDF+;[2
DSC#SC
RNRPs25[RR:=';j'
MSC8VRH;R
RCRM8DbFF;R
RskC0sPMRN
s;CRM8b;N8
MVkOF0HMCRo0H_I8_0EUH5I8:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=I0H8E;/U
HRRV5R5I0H8EFRl82RURc>R2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCI0_HE80_
U;VOkM0MHFR0oC_8IH0.E_58IH0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:I=RHE80/
.;RCRs0MksRDPN;M
C8CRo0H_I8_0E.V;
k0MOHRFMo_C0I0H8EH5I8R0E:MRH0CCoss2RCs0kMCRDVP0FC0s__H.R#N
PsLHNDPCRN:DRRVDC0CFPs__0.L;
CMoH
PRRN4D52=R:R0oC_8IH0.E_58IH0;E2
HRRVIR5HE80R8lFR=.RRRj20MEC
RRRRDPN5Rj2:j=R;R
RCCD#
RRRRDPN5Rj2:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0H_I8;0E
MVkOF0HMCRo0H_I850EI0H8ERR:HCM0o2CsR0sCkRsMD0CVFsPC_H0R#N
PsLHNDPCRN:DRRVDC0CFPsR_0:5=Rjj,R,,RjR;j2
oLCHRM
RDPN5Rd2:o=RCI0_HE80_IU5HE802R;
R#ONCIR5HE80R8lFRRU2HR#
RCIEMRRc|RRd=P>RN.D52=R:R
4;RERIC.MRRR=>P5ND4:2R=;R4
IRRERCM4>R=RDPN5Rj2:4=R;R
RIMECREF0CRs#=M>Rk;DD
CRRMO8RN;#C
sRRCs0kMNRPDC;
Mo8RCI0_HE80;F
OMN#0M#0R_8IH0NE_s$sNRD:RCFV0P_Cs0=R:R0oC_8IH0IE5HE802O;
F0M#NRM0#H_I8_0ENNss$c_nRD:RCFV0P_Cs0R_.:o=RCI0_HE8058IH0;E2
MVkOF0HMCRo0k_Ml._4UC58b:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=80CbE./4UR;
RRHV5C58bR0ElRF842.UR4>R4R.20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_U4.;k
VMHO0FoMRCD0_CFV0P_Csn8c5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#C
Lo
HMRCRs0Mks5b8C0lERF48R.;U2
8CMR0oC_VDC0CFPsc_n;k
VMHO0FoMRCM0_knl_cC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=R4N.RM88RCEb0Rc>RU02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC5b8C0:ERR0HMCsoC;NRlGRR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbERR-lRNG>j=R2ER0CRM
RPRRN:DR=CR8bR0E-NRlGR;
R#CDCR
RRNRPD=R:Rb8C0
E;RMRC8VRH;R
RskC0sPM5N;D2
8CMR0oC_VDC0CFPsV;
k0MOHRFMo_C0M_kld8.5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=cNURM88RCEb0R4>Rn02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_kdl_.V;
k0MOHRFMo_C0M_kl48n5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4NnRM88RCEb0Rj>R2ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Mln_4;-
-O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5855CEb0R4-R2RR/dR.2+5R55b8C0-ERRR42lRF8dR.2/nR42R2;R-R-RFyRVqR)vXd.4O1RC#DDRCMC8RC8
MOF#M0N0kRMlC_OD4D_.:URR0HMCsoCRR:=o_C0M_kl45.U80CbE
2;O#FM00NMRVDC0CFPsc_nRH:RMo0CC:sR=CRo0C_DVP0FCns_cC58b20E;F
OMN#0MM0RkOl_C_DDn:cRR0HMCsoCRR:=o_C0M_klnDc5CFV0P_Csn;c2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,ncR2nc;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bC4R.UHN#Rs$sNRk5MlC_OD4D_.8URF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bnC_c#RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdH.R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_R4nHN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k4#_.:URR0Fk_#Lk_b0$C._4UR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kn#_cRR:F_k0L_k#0C$b_;ncRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_k4#_nRR:F_k0L_k#0C$b_;4nRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNRF#_kC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD._4UFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CLMNDRC#VRFs0-sH#00NC##
HNoMDkRF0M_C_Rnc:0R#8F_Do;HO
o#HMRNDF_k0CdM_.RR:#_08DHFoO#;
HNoMDkRF0M_C_R4n:0R#8F_Do;HO
o#HMRND#s_I0M_CR#:R0D8_FOoH_OPC05FsM_klODCD_U4.RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rnc:0R#8F_Do;HO
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRND#M_H_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNRF#_ks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD_R#Ns8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#CqsR7
7)#MHoNDDRFNI_8R8s:0R#8F_Do_HOP0COFns5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82O#FM00NMRLD#_8IH0:ERR0HMCsoCRR:=I0H8E*-U5I#_HE80_sNsNd$522-4-#c*_8IH0NE_s$sN5-.2._*#I0H8Es_Ns5N$4#2-_8IH0NE_s$sN5;j2
b0$ClR0bs_NsUN$RRH#NNss$#R5_8IH0NE_s$sN5-d24FR8IFM0RRj2F#VR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
o#HMRND0_lbU._d,lR0b__U4:nRRb0l_sNsN;$U
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
RR
RzRcd:VRHR85N8ss_CRo2oCCMsCN0RR--oCCMsCN0RFLDOs	RNRl
R-RR-VRQR8N8s8IH0<ERRFOEH_OCI0H8E#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8R8s<"=Rjjjjjjjjjjjjj&"RR7q7)25j;R
RRRRRRFRDIN_I8R8s<"=Rjjjjjjjjjjjjj&"RR_N8s5Coj
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjjjjjj&"RR7q7)R548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjjjjj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjjjjjj&"RR7q7)R5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjjjjj"RR&Ns8_C.o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjj"jjRq&R757)dFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjj"jjRq&R757)cFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjjjjjj&"RR7q7)R568MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjjj&"RR_N8s5Co6FR8IFM0R;j2
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRNs88I0H8ERR=(o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjjjjj&"RR7q7)R5n8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjjjjjj"RR&Ns8_Cno5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjjj"jjRq&R757)(FR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjjj&"RR_N8s5Co(FR8IFM0R;j2
RRRR8CMRMoCC0sNC(Rz;R
RRURzRRR:H5VRNs88I0H8ERR=go2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj"jjRq&R757)UFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=jR"jjjj"RR&Ns8_CUo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zU
RRRRRzgRH:RVNR58I8sHE80R4=Rjo2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jjRj"&7Rq7g)5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<Rj"jjRj"&8RN_osC58gRF0IMF2Rj;R
RRMRC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<="jjj"RR&q)775R4j8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
RRRR8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0RC
RRRRRDRRFsI_Ns88RR<=""jjRq&R757)484RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&8RN_osC5R448MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;44
RRRR.z4RRR:H5VRNs88I0H8ERR=4Rd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR''RR&q)775R4.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&8RN_osC5R4.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RRR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=7Rq74)5dFR8IFM0R;j2
RRRRRRRRIDF_8IN8<sR=8RN_osC5R4d8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRR8CMRMoCC0sNC4Rz6
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C)sR_z7ma#RkHRMo)B_mpRi
RzRR4RnR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s4Co2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s4Co;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRR(z4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C;o4
RRRR8CMRMoCC0sNC4Rz(
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7V)RFIsRsCH0RHk#MBoRpRi
RzRR4RUIRH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4RzU
I;RRRRzI4gRH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR8RN_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4;gI
R
RR-R-R0 GsDNRFOoHRsVFRN7kDFRbsO0RN
#CSR--7MFRFM0RCRC80#EHRsVFRRMFokDFCFRDoRHOO8FMHF0HM-
-RRRRzosCRb:RsCFO#B#5pRi2LHCoM-
-RRRRRVRHRp5Bie'  RhaNRM8BRpi=4R''02RE
CM-R-RRRRRRh7Q_b0lRR<=7;Qh
R--RRRRRqR)7_7)0Rlb<q=R7;7)
R--RRRRRqRW7_7)0Rlb<N=R8C_so-;
-RRRRRRRW0 _l<bR= RW;-
-RRRRRMRC8VRH;-
-RRRRCRM8bOsFC;##
R
RRlRzk:GRRFbsO#C#50Fk_osC2R
RRRRRLHCoM-
-RRRRRRRRH5VRW7q7)l_0bRR=)7q7)l_0bMRN8 RW_b0lR'=R4R'20MEC
R--RRRRRRRRR0Fk_osC4=R<Rh7Q_b0l;-
-RRRRRRRRCCD#
RRRRRRRRFRRks0_CRo4<F=Rks0_CIo5HE80-84RF0IMF2Rj;-
-RRRRRRRRCRM8H
V;RRRRCRM8bOsFC;##
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n114_4R
RR4RzURR:H5VROHEFOIC_HE80R4=R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RRRRRORzE:	RRRHV58RN8HsI8R0E>cR42CRoMNCs0RC
RRRRRRRRRkRRO:D	RFbsO#C#5iBp2R
RRRRRRRRRRLRRCMoH
RRRRRRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRRRRR8sN8ss_CNo58I8sHE80-84RF0IMFcR42=R<R7q7)85N8HsI8-0E4FR8IFM0R24c;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8bOsFC;##
RSSR8CMRMoCC0sNCORzE
	;RRRRRRRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjz.RH:RVNR58I8sHE80R4>Rco2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns88_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
j;RRRR-Q-RVNR58I8sHE80RR<=4Rc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4z.;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRR.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vn_4dXUc4:7RRv)qA_4n114_4R
RRRRRRRRRRRRRRFRbsl0RN5bR75Qqj=2R>MRH_osC5,[2R7q7)=qR>FRDIN_I858s48dRF0IMF2Rj,QR7A>R=R""j,7Rq7R)A=D>RFsI_Ns885R4d8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25jRR=>F_k0L4k#5[H,2
2;
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
.;RRRRRRRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1.1R.
RzRR.:dRRRHV5FOEH_OCI0H8ERR=.o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRRORzER	:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRRRRRDkO	b:RsCFO#B#5p
i2RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRRRRRsRRNs88_osC58N8s8IH04E-RI8FMR0F4Rd2<q=R757)Ns88I0H8ER-48MFI04FRd
2;RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRMRC8sRbF#OC#S;
SMRC8CRoMNCs0zCRO;E	
RRRRRRRRcz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRRRRR.Rz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8N8sC_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.6
RRRRR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRRRRRR.RznRR:H5VRNs88I0H8E=R<R24dRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRRRRR8CMRMoCC0sNC.RznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRRRRRzR.(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAqUv_4Xg..:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)v4_Ug..X7RR:)Aqv41n_.._1
RRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A254RR=>F_k0L.k#5.H,*4[+27,RmjA52>R=R0Fk_#Lk.,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co.2*[RR<=F_k0L.k#5.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[.*+R42<F=RkL0_k5#.H*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
(;RRRRRRRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RR

RRRRR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1c1Rc
RzRR.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRRzRRO:E	RRHV58N8s8IH0>ERR24.RMoCC0sNCR
RRRRRRRRRRORkDR	:bOsFC5##B2pi
RRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRRRRRs8N8sC_so85N8HsI8-0E4FR8IFM0R24.RR<=q)7758N8s8IH04E-RI8FMR0F4;.2
RRRRRRRRRRRRCRRMH8RVR;
RRRRRRRRRCRRMb8RsCFO#
#;SRSRCRM8oCCMsCN0REzO	R;
RRRRRzRR.:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERR24.RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRRRRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRN5s8_8ss5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRR8CMRMoCC0sNCdRzjR;
R-RR-VRQR85N8HsI8R0E<4=R.M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRRRRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;d4
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRRRRRdRz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRARR)_qvcnjgXRc7:qR)vnA4__1c1Rc
RRRRRRRRRRRRRbRRFRs0lRNb5q7QRR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7R)q=D>RFII_Ns885R448MFI0jFR27,RQ=AR>jR"j"jj,7Rq7R)A=D>RFsI_Ns885R448MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25dRR=>F_k0Lck#5RH,c+*[dR2,75mA.=2R>kRF0k_L#Hc5,[c*+,.2RR
RRRRRRRRRRRRRRmR7A254RR=>F_k0Lck#5cH,*4[+27,RmjA52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';
RRRRRRRRRRRR8CMRMoCC0sNCdRz.R;
RRRRRCRRMo8RCsMCNR0Cz;.g
RRRR8CMRMoCC0sNC.RzU
;
RRRRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1_
1gRRRRzRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRRRRRz	OE:VRHR85N8HsI8R0E>4R42CRoMNCs0RC
RRRRRRRRRkRRO:D	RFbsO#C#5iBp2R
RRRRRRRRRRLRRCMoH
RRRRRRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRRRRR8sN8ss_CNo58I8sHE80-84RF0IMF4R42=R<R7q7)85N8HsI8-0E4FR8IFM0R244;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8bOsFC;##
RSSR8CMRMoCC0sNCORzE
	;RRRRRRRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>4R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRR6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns88_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
6;RRRR-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRRnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rnzd;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRRd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRAv)q_c.jU7XUR):Rq4vAng_1_
1gRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5g[R+(8MFI0gFR*,[2R7q7)=qR>FRDIN_I858s48jRF0IMF2Rj,QR7A>R=Rj"jjjjjj,j"R7q7)=AR>FRDIN_s858s48jRF0IMF2Rj,R
RRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A25(RR=>F_k0LUk#5UH,*([+27,RmnA52>R=R0Fk_#LkU,5HU+*[nR2,
RRRRRRRRRRRRRRRRA7m5R62=F>RkL0_k5#UH*,U[2+6,mR7A25cRR=>F_k0LUk#5UH,*c[+27,RmdA52>R=R0Fk_#LkU,5HU+*[dR2,
RRRRRRRRRRRRRRRRA7m5R.2=F>RkL0_k5#UH*,U[2+.,mR7A254RR=>F_k0LUk#5UH,*4[+27,RmjA52>R=R0Fk_#LkU,5HU2*[,R
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7ujq52>R=R_HMs5Cog+*[UR2,7AQuRR=>",j"Ru7mq>R=RCFbM7,Rm5uAj=2R>NRbs$H0_#LkU,5HR2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRMRC8CRoMNCs0zCRd
(;RRRRRRRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RRRRRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_41U_4RU
RzRRd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRRRRRz	OE:VRHR85N8HsI8R0E>jR42CRoMNCs0RC
RRRRRRRRRkRRO:D	RFbsO#C#5iBp2R
RRRRRRRRRRLRRCMoH
RRRRRRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRRRRR8sN8ss_CNo58I8sHE80-84RF0IMFjR42=R<R7q7)85N8HsI8-0E4FR8IFM0R24j;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRCRM8bOsFC;##
RSSR8CMRMoCC0sNCORzE
	;RRRRRRRRzRdg:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>jR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRRRRRjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns88_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRMRC8CRoMNCs0zCRc
j;RRRR-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRRRRR4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0R4zc;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRRRRRzRRc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXn:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRRRRRqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2R,
RRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRR
RRRRRRRRRRRRRRmR7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RR
RRRRRRRRRRRRRRmR7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RR
RRRRRRRRRRRRRRmR7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RR
RRRRRRRRRRRRRRmR7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RRRRRRRRRRRRRRRRR75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RR
RRRRRRRRRRRRRRmR7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mq>R=RCFbM7,Rm5uA4=2R>NRbs$H0_#Lk4Hn5,*R.[2+4,mR7ujA52>R=RsbNH_0$L4k#n,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co4[U*2=R<R0Fk_#Lk4Hn5,*4n[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R42<F=RkL0_kn#454H,n+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R.2<F=RkL0_kn#454H,n+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rd2<F=RkL0_kn#454H,n+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rc2<F=RkL0_kn#454H,n+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R62<F=RkL0_kn#454H,n+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rn2<F=RkL0_kn#454H,n+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R(2<F=RkL0_kn#454H,n+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+RU2<F=RkL0_kn#454H,n+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rg2<F=RkL0_kn#454H,n+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24jRR<=F_k0L4k#n,5H4[n*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+4<2R=kRF0k_L#54nHn,4*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24.RR<=F_k0L4k#n,5H4[n*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+d<2R=kRF0k_L#54nHn,4*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24cRR<=F_k0L4k#n,5H4[n*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+6<2R=kRF0k_L#54nHn,4*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24nRR<=bHNs0L$_kn#45.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[(+42=R<RsbNH_0$L4k#n,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.zc;R
RRRRRRMRC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nd_1nz
SdRUN:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SRRRRREzO	H:RVNR58I8sHE80Rg>R2CRoMNCs0SC
SRRRRDkO	b:RsCFO#B#5p
i2SRSSLHCoMS
SSHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
SSSRRRRs8N8sC_so85N8HsI8-0E4FR8IFM0RRg2<q=R757)Ns88I0H8ER-48MFI0gFR2S;
SRSRCRM8H
V;SCSSMb8RsCFO#
#;SRSRCRM8oCCMsCN0REzO	S;
RRRRzNdgRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SSjzcNRR:H5VRNs88I0H8ERR>go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRSSRFRRkC0_M25HRR<='R4'IMECRN5s8_8ss5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc;jN
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SS4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0CzNc4;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSScR.N:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
SSSSqA)v4_6..Xd7RR:)Aqv41n_d1n_dRn
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7q7)RR=>D_FII8N8sR5U8MFI0jFR2
,RSSSS7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSSq7mRR=>FMbC,mR7A45d2>R=R0Fk_#LkdH.5,*d.[4+d27,RmdA5j=2R>kRF0k_L#5d.H.,d*d[+j
2,SSSS75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2S,
S7SSm.A5n=2R>kRF0k_L#5d.H.,d*.[+nR2,75mA.R62=F>RkL0_k.#d5dH,.+*[.,62RA7m52.cRR=>F_k0Ldk#.,5Hd[.*+2.c,S
SSmS7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
SSSSA7m52.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7Ag542>R=R0Fk_#LkdH.5,*d.[g+427,Rm4A5U=2R>kRF0k_L#5d.H.,d*4[+U
2,SSSS75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42S,
S7SSm4A5c=2R>kRF0k_L#5d.H.,d*4[+cR2,75mA4Rd2=F>RkL0_k.#d5dH,.+*[4,d2RA7m524.RR=>F_k0Ldk#.,5Hd[.*+24.,SR
S7SSm4A54=2R>kRF0k_L#5d.H.,d*4[+4R2,75mA4Rj2=F>RkL0_k.#d5dH,.+*[4,j2RA7m5Rg2=F>RkL0_k.#d5dH,.+*[gR2,
SSSSA7m5RU2=F>RkL0_k.#d5dH,.+*[UR2,75mA(=2R>kRF0k_L#5d.H.,d*([+27,RmnA52>R=R0Fk_#LkdH.5,*d.[2+n,SR
S7SSm6A52>R=R0Fk_#LkdH.5,*d.[2+6,mR7A25cRR=>F_k0Ldk#.,5Hd[.*+,c2RA7m5Rd2=F>RkL0_k.#d5dH,.+*[dR2,
SSSSA7m5R.2=F>RkL0_k.#d5dH,.+*[.R2,75mA4=2R>kRF0k_L#5d.H.,d*4[+27,RmjA52>R=R0Fk_#LkdH.5,*d.[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq>R=R_HMs5Cod[n*+Rd68MFI0dFRn+*[d,.2Ru7QA>R=Rj"jj,j"Ru7mq>R=RCFbM7,Rm5uAd=2R>NRbs$H0_#LkdH.5,[c*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA25.RR=>bHNs0L$_k.#d5cH,*.[+27,Rm5uA4=2R>NRbs$H0_#LkdH.5,[c*+,42Ru7mA25jRR=>bHNs0L$_k.#d5cH,*2[2;R
RRRRRRRRRRRRRRkRF0C_son5d*R[2<F=RkL0_k.#d5dH,.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+2=R<R0Fk_#LkdH.5,*d.[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*c[+2=R<R0Fk_#LkdH.5,*d.[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*n[+2=R<R0Fk_#LkdH.5,*d.[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*U[+2=R<R0Fk_#LkdH.5,*d.[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+j<2R=kRF0k_L#5d.H.,d*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+.<2R=kRF0k_L#5d.H.,d*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+c<2R=kRF0k_L#5d.H.,d*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+n<2R=kRF0k_L#5d.H.,d*4[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*4[+U<2R=kRF0k_L#5d.H.,d*4[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+j<2R=kRF0k_L#5d.H.,d*.[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+.<2R=kRF0k_L#5d.H.,d*.[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+c<2R=kRF0k_L#5d.H.,d*.[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+n<2R=kRF0k_L#5d.H.,d*.[+nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*.[+U<2R=kRF0k_L#5d.H.,d*.[+UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+j<2R=kRF0k_L#5d.H.,d*d[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+.<2R=NRbs$H0_#LkdH.5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_son5d*d[+c<2R=NRbs$H0_#LkdH.5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0R.zcNR;
RRRRRCRRMo8RCsMCNR0CzNdg;R
RRMRC8CRoMNCs0zCRd;UN
CRRMo8RCsMCNR0Cz;cd
zRRcRc:H5VRMRF0Ns88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<(#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jjjjj&"RRN#_8C_so25j;R
RRMRC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8N8s=R<Rj"jj"jjR#&R__N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj&"RRN#_8C_soR5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jRj"&_R#Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
cSzSH:RVNR58I8sHE80R6=R2CRoMNCs0SC
SIDF_8N8s=R<Rj"j"RR&#8_N_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;SSz6:VRHR85N8HsI8R0E=2RnRMoCC0sNCS
SD_FINs88RR<='Rj'&_R#Ns8_C6o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<#=R__N8s5ConFR8IFM0R;j2
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR(RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRRH#_MC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRR#M_H_osCRR<=7;Qh
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRzgRH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=#k_F0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<#=R_0Fk_osC;R
RRMRC8CRoMNCs0zCR4
j;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBiR
RR4Rz4:RRRRHV58N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRR#8_N_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz4R;
RzRR4:.RRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRR#8_N_osCRR<=q)77;R
RRMRC8CRoMNCs0zCR4
.;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4d:FRVsRRHH5MRM_klODCD_U4.R4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRcz4RH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRR#RR_0Fk_5CMH<2R=4R''ERIC5MR#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRR_R#I_s0CHM52=R<RRW IMECR_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rcz4;R
RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4Rz6RR:H5VRNs88I0H8E=R<RR(2oCCMsCN0
RRRRRRRRRRRRRRRRF#_kC0_M25HRR<=';4'
RRRRRRRRRRRRRRRRI#_sC0_M25HRR<=W
 ;RRRRRRRRCRM8oCCMsCN0R6z4;R
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRzRR4:nRRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qv.:URRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*.RU2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H442*.RU,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.v4URR:Xv)q4X.U4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5Co[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6R2,q=nR>FRDI8_N8ns52S,
SSSSSWRR >R=RI#_sC0_M25H,BRWp=iR>pRBim,RRR=>F_k0L_k#45.UH2,[2R;
RRRRRRRRRRRRR#RR_0Fk_osC5R[2<F=RkL0_k4#_.HU5,R[2IMECR_5#F_k0CHM52RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRRMRC8CRoMNCs0zCR4Rd;RRRRRRRRR
RRRRRRRRR
R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR(z4RH:RVMR5kOl_C_DDn=cRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>(M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4RzU:NRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mc_nRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4NR;
RRRRRzRR4RUL:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_U4.Rj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECR#55__N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5#8_N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UL
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRgz4RH:RVNR58I8sHE80RR<=no2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CnM_c=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rnc<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;4g
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_.:VRHR_5#I0H8Es_Ns_N$n4c52RR>jo2RCsMCN
0CRRRRRRRRzR.j:FRVsRR[H5MR#H_I8_0ENNss$c_n5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RzqcvnRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U42.UR"&RW&"RR0HMCsoC'NHloIC5HE80R.-R*-[RRR.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERR[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR.1
RRRRRRRRRRRRRRRRsbF0NRlb7R54>R=RH#_MC_soH5I8-0E.-*[4R2,7=jR>_R#HsM_CIo5HE80-[.*-,.2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c,6RqRR=>D_FINs885,62
SSSSRSSRRW =I>RsC0_Mc_n,BRWp=iR>pRBim,R4>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-4,jRmRR=>F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-2.2;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-.[2-4RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-[.*-R.2<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[.I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNC.RzjS;
SMRC8CRoMNCs0zCRO_E	.S;
SORzE4	_RH:RV#R5_8IH0NE_s$sN_5ncj>2RRRj2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERR#.*_8IH0NE_s$sN_5nc4-2RRR42& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.Rn+Rc8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERR#.*_8IH0NE_s$sN_5nc4;22
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_soH5I8-0E._*#I0H8Es_Ns_N$n4c522-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,S
SSSSSR RWRR=>I_s0CnM_cW,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.#H_I8_0ENNss$c_n5-424;22
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#.*_8IH0NE_s$sN_5nc442-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.#H_I8_0ENNss$c_n5-424I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNCORzE4	_;R
SRRRRCRM8oCCMsCN0R(z4;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:4RRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN..RH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.N
RRRRRRRR.z.LRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_c=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M._dRR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z.LR;
RRRRRzRR.R.O:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
O;RRRRRRRRz8..RH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCDc_nRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDc_n2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F6=2RRlMk_DOCDc_n2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
8;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.d:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RW;R
RRRRRRMRC8CRoMNCs0zCR.
d;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:URRRHV5I#_HE80_sNsNd$52RR>jo2RCsMCN
0CSOSzED	_C:6RRRHV58IH0>ER=*RU#H_I8_0ENNss$25dR8NMR8IH0>ER=2RURMoCC0sNCR
RRRRRRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR+U
2;RRRRRRRRRRRRRRRRRRRRLHCoMS
SRRRRzv)qd:.RRqX)vXd.US1
SRSRRFRbsl0RN5bR7>R=R8bN5H#_MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.HR[2<0=RlUb__5d.jH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R[-R*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-[R5-*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_soH5I8-0ED_#LI0H8E*-U[R+(8MFI0IFRHE80-LD#_8IH0UE-*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=Rb0l_dU_.25[2S;
SRSRR#RN#MHoRV:RFHsR[MRHR8(RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.H,I8-0ED_#LI0H8E*-U[[+H2=R<Rb0l_dU_.25[52H[;R
RRRRRRRRRRRRRRRRR#k_F0C_soH5I8-0ED_#LI0H8E*-U[[+H2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E#-DLH_I8-0EU+*[HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	D;C6
zSSO_E	oR06:VRHRH5I8R0E>U=RR8NMR8IH0lERFU8RRR>=6o2RCsMCN
0CRRRRRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbU._d5I#_HE80_sNsNd$522-42S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Ud#.5_8IH0NE_s$sN5-d24H25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRzR.U:FRVsRR[H#MR_8IH0NE_s$sN5-d2.FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C5*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC[55+*42U
2;RRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRR)Rzq.vdRX:R)dqv.1XURR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RH#_MC_so*5U[R+(8MFI0UFR*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=Rb0l_dU_.25[2S;
SNSS#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdU.,*H[+[<2R=lR0b__Ud[.52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CUo5*H[+[<2R=kRF0k_L#._d5lMk_DOCD._d,[U*+2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHloUC52R;
RRRRRRRRRRRRRRRRRLRRCMoH
RSSRzRR)dqv.RR:Xv)qdU.X1S
SSRRRRsbF0NRlb7R5RR=>b5N8#M_H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_.25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#._d5lMk_DOCD._d,2H[RR<=0_lbU._d55j2H;[2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
CSSMo8RCsMCNR0Cz	OE_
M;SMSC8CRoMNCs0zCRO_E	US;
SEzO	R_c:VRHR_5#I0H8Es_Ns5N$.>2RRRj2oCCMsCN0
RRRRRRRRcz._:cRRRHV58IH0>ER=2RcRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>_R#HsM_Cdo527,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,
SSSSRSSRRmd=F>RkL0_kd#_.k5MlC_ODdD_.2,d,.RmRR=>F_k0L_k#dM.5kOl_C_DDd..,2S,
SSSSSmRR4>R=R0Fk_#Lk_5d.M_klODCD_,d.4R2,m=jR>kRF0k_L#._d5lMk_DOCD._d,2j2;R
RRRRRRRRRRRRRR_R#F_k0s5Cod<2R=kRF0k_L#._d5lMk_DOCD._d,Rd2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_5d.M_klODCD_,d..I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_kd#_.k5MlC_ODdD_.2,jRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.cc_;R
RRRRRR.RzcR_d:VRHRH5I8R0E=2RdRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRd.:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzq.vdRX:R)dqv.1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>jR''7,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,
SSSSRSSRRmd=F>Rb,CMRRm.=F>RkL0_kd#_.k5MlC_ODdD_.2,.,S
SSSSSR4RmRR=>F_k0L_k#dM.5kOl_C_DDd4.,2m,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRRF#_ks0_C.o52=R<R0Fk_#Lk_5d.M_klODCD_,d..I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so254RR<=F_k0L_k#dM.5kOl_C_DDd4.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rj2<F=RkL0_kd#_.k5MlC_ODdD_.2,jRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.dc_;S
SCRM8oCCMsCN0REzO	;_c
zSSO_E	.RR:H5VR#H_I8_0ENNss$254Rj>R2CRoMNCs0RC
RRRRRzRR.:cRRsVFRH[RM#R5_8IH0NE_s$sN5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNCH5I8-0EU_*#I0H8Es_Ns5N$d.2-*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:)dqv.1X.RR
RRRRRRRRRRRRRRFRbsl0RN5bR7=jR>_R#HsM_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.R2,7=4R>_R#HsM_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[4R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,Rj>R=R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.H,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2
2;RRRRRRRRRRRRRRRR#k_F0C_soH5I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-U#H_I8_0ENNss$25d-[.*-R42IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_CIo5HE80-#U*_8IH0NE_s$sN5-d2.-*[.<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*I#_HE80_sNsNd$52*-.[2-.RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
c;SMSC8CRoMNCs0zCRO_E	.S;
SEzO	R_4:VRHR_5#I0H8Es_Ns5N$j>2RRRj2oCCMsCN0
RRRRRRRRcz.RH:RVIR5HE80R8lFR=URRR42oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRR,d.Rb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:qR)vXd.4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CojR2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBim,RRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
4;RRRRCRM8oCCMsCN0R4z.;RRRRRRRR
RR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR.:6RRRHV5lMk_DOCDn_4R4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nN
RRRRRRRRnz.LRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58R#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=jR''N2RM58R#8_N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL.n;R
RRRRRR.Rzn:ORRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRNjRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85N#_8C_so25nR'=RjR'2NRM85N#_8C_so256R'=R4R'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.OR;
RRRRRzRR.Rn8:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR_5#Ns8_Cno52RR='2j'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8#R5__N8s5Con=2RR''j2MRN8#R5__N8s5Co6=2RR''j2MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
8;RRRRRRRRzC.nRH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECR#55__N8s5Con=2RR''42MRN8#R5__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC5Rn2=4R''N2RM58R#8_N_osC5R62=4R''N2RMR8R5N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzC.n;R
RRRRRR.Rzn:VRRRHV58N8s8IH0=ERRN(RMM8RkOl_C_DDn=cRRN4RMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5N#_8C_so25nR'=R4R'2NRM85N#_8C_so256R'=RjR'2NRM85N#_8C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5_5#Ns8_Cno52RR='24'R8NMR_5#Ns8_C6o52RR='2j'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.VR;
RRRRRzRR.Rno:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=RRjNRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5_5#Ns8_C6o52RR='24'R8NMR_5#Ns8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECR#55__N8s5Co6=2RR''42MRN8#R5__N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
o;RRRRRRRRzE.nRH:RVNR58I8sHE80R6=RR8NMRlMk_DOCD._dRR/=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5#8_N_osC58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
E;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.(:VRHR85N8HsI8R0E<c=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<=';4'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RW;R
RRRRRRMRC8CRoMNCs0zCR.
(;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00SC
RRRRz	OE_:URRRHV5I#_HE80_sNsNd$52RR>jo2RCsMCN
0CSOSzED	_C:6RRRHV58IH0>ER=*RU#H_I8_0ENNss$25dR8NMR8IH0>ER=2RURMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Hn,[<2R=lR0b__U4jn52[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRRF#_ks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RM_R#I0H8Es_Ns5N$d42-RI8FMR0F4CRoMNCs0RC
RRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R[-R*RU2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80R5-R[2-4*;U2
RRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRRzRR)4qvnRR:Xv)q4UnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>_R#HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,RRm=0>RlUb__54n[;22
SSSRRRRNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nI0H8E#-DLH_I8-0EU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoI0H8E#-DLH_I8-0EU+*[HR[2<F=RkL0_k4#_nk5MlC_OD4D_nH,I8-0ED_#LI0H8E*-U[[+H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRCRRMo8RCsMCNR0CNH##o
M;RRRRRRRRRRRRCRM8oCCMsCN0RUz.;S
SCRM8oCCMsCN0REzO	C_D6S;
SEzO	0_o6RR:H5VRI0H8E=R>RNURMI8RHE80R8lFR>UR=2R6RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E+2RU;R
RRRRRRRRRRCRLo
HMSRSRR)Rzqnv4RX:R)4qvn1XU
SSSRRRRb0FsRblNRR57=b>RN#85__HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n_5#I0H8Es_Ns5N$d42-2
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54n#H_I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRR#RR_0Fk_osC52H[RR<=F_k0L_k#4Mn5kOl_C_DD4Hn,[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHM#H_I8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5U[*2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vR4n:)RXqnv4XRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>#M_H_osC5[U*+8(RF0IMF*RU[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=Rb0l_4U_n25[2S;
SNSS#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4Un,*H[+[<2R=lR0b__U4[n52[5H2R;
RRRRRRRRRRRRRRRRRF#_ks0_CUo5*H[+[<2R=kRF0k_L#n_45lMk_DOCDn_4,[U*+2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRMRC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRCRRMo8RCsMCNR0Cz;.U
CSSMo8RCsMCNR0Cz	OE_6o0;S
Sz	OE_:MRRRHV58IH0<ERRRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vR4n:)RXqnv4X
U1SRSSRbRRFRs0lRNb5=7R>NRb8_5#HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbUn_452j2;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54njH25[
2;RRRRRRRRRRRRRRRRR_R#F_k0s5CoHR[2<F=RkL0_k4#_nk5MlC_OD4D_n[,H2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;SMSC8CRoMNCs0zCRO_E	MS;
S8CMRMoCC0sNCORzEU	_;S
Sz	OE_:cRRRHV5I#_HE80_sNsN.$52RR>jo2RCsMCN
0CRRRRRRRRz_.gcRR:H5VRI0H8E=R>RRc2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHlojC52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)4qvnRR:)4qvn1XcRR
RRRRRRRRRRRRRRFRbsl0RN5bR7=dR>_R#HsM_Cdo527,R.>R=RH#_MC_so25.,4R7RR=>#M_H_osC5,42RR7j=#>R__HMs5Coj
2,SRSSRRRRRRRRRRRRRRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRS
SSSSSRdRmRR=>F_k0L_k#4Mn5kOl_C_DD4dn,2m,R.>R=R0Fk_#Lk_54nM_klODCD_,4n.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,,42RRmj=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRR#RR_0Fk_osC5Rd2<F=RkL0_k4#_nk5MlC_OD4D_n2,dRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Co.<2R=kRF0k_L#n_45lMk_DOCDn_4,R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRF#_ks0_C4o52=R<R0Fk_#Lk_54nM_klODCD_,4n4I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRR#k_F0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.gcR;
RRRRRzRR.dg_RH:RVIR5HE80Rd=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlocC52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4nc
1RRRRRRRRRRRRRRRRRb0FsRblNRd57RR=>',j'RR7.=#>R__HMs5Co.R2,7=4R>_R#HsM_C4o527,Rj>R=RH#_MC_so25j,S
SSRRRRRRRRRRRRqRRj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi
,RSSSSSRSRm=dR>bRFCRM,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRR#k_F0C_so25.RR<=F_k0L_k#4Mn5kOl_C_DD4.n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC5R42<F=RkL0_k4#_nk5MlC_OD4D_n2,4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRR_R#F_k0s5Coj<2R=kRF0k_L#n_45lMk_DOCDn_4,Rj2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC.Rzg;_d
CSSMo8RCsMCNR0Cz	OE_
c;SOSzE.	_RH:RV#R5_8IH0NE_s$sN5R42>2RjRMoCC0sNCR
RRRRRRdRzjRR:VRFs[MRHR_5#I0H8Es_Ns5N$4-2RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8E*-U#H_I8_0ENNss$25d-[.*-R.2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80-#U*_8IH0NE_s$sN5-d2.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4.nX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,.2RR74=#>R__HMs5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-,42RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piRRmj=F>RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*.[-2S,
SSSSSmRR4>R=R0Fk_#Lk_54nM_klODCD_,4nI0H8E*-U#H_I8_0ENNss$25d-[.*-242;R
RRRRRRRRRRRRRR_R#F_k0s5CoI0H8E*-U#H_I8_0ENNss$25d-[.*-R42<F=RkL0_k4#_nk5MlC_OD4D_nH,I8-0EU_*#I0H8Es_Ns5N$d.2-*4[-2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRR#RR_0Fk_osC58IH0UE-*I#_HE80_sNsNd$52*-.[2-.RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-#U*_8IH0NE_s$sN5-d2.-*[.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rjzd;S
SCRM8oCCMsCN0REzO	;_.
zSSO_E	4RR:H5VR#H_I8_0ENNss$25jRj>R2CRoMNCs0RC
RRRRRzRRd:4RRRHV58IH0lERFU8RR4=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo4C52R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=#>R__HMs5CojR2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,m>R=R0Fk_#Lk_54nM_klODCD_,4nj;22
RRRRRRRRRRRRRRRRF#_ks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R4zd;S
SCRM8oCCMsCN0REzO	;_4
RRRRMRC8CRoMNCs0zCR.R6;RRRRRRRRRR
RR8CMRMoCC0sNCcRzcC;
MN8RsHOE00COkRsCMsF_IE_OC;O	
-
-

------R#pN0lRHblDCCNM00MHFRRH#8NCVk
D0-N-
sHOE00COkRsC#CCDOs0_NFlRVqR)vW_)R
H#ObFlFMMC0)RXq.v4U1X4
FRbs50R
RRRmRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRRq:6RRRHM#_08DHFoOR;
RnRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;


ObFlFMMC0)RXqcvnX
.1RsbF0
R5RmRRjRR:FRk0#_08DHFoOR;
R4RmRF:Rk#0R0D8_FOoH;R
RRRqj:MRHR8#0_oDFH
O;RqRR4RR:H#MR0D8_FOoH;R
RRRq.:MRHR8#0_oDFH
O;RqRRdRR:H#MR0D8_FOoH;R
RRRqc:MRHR8#0_oDFH
O;RqRR6RR:H#MR0D8_FOoH;R
RRR7j:MRHR8#0_oDFH
O;R7RR4RR:H#MR0D8_FOoH;R
RRpWBiRR:H#MR0D8_FOoH;R
RRRW :MRHR8#0_oDFHRO
2C;
MO8RFFlbM0CM;O

FFlbM0CMRqX)vXd.cR1
b0FsRR5
RjRmRF:Rk#0R0D8_FOoH;R
RRRm4:kRF00R#8F_Do;HO
RRRm:.RR0FkR8#0_oDFH
O;RmRRdRR:FRk0#_08DHFoOR;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7:jRRRHM#_08DHFoOR;
R4R7RH:RM0R#8F_Do;HO
RRR7:.RRRHM#_08DHFoOR;
RdR7RH:RM0R#8F_Do;HO
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
lOFbCFMMX0R)dqv.1XU
b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RcRqRH:RM0R#8F_Do;HO
RRR7RR:H#MR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
RRRWiBpRH:RM0R#8F_Do;HO
RRRW: RRRHM#_08DHFoO2
R;M
C8FROlMbFC;M0
F
OlMbFCRM0Xv)q4UnX1b
RFRs05R
RR:mRR0FkR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RjRqRH:RM0R#8F_Do;HO
RRRq:4RRRHM#_08DHFoOR;
R.RqRH:RM0R#8F_Do;HO
RRRq:dRRRHM#_08DHFoOR;
RRR7:MRHR8#0_oDFHPO_CFO0sR5(8MFI0jFR2R;
RBRWp:iRRRHM#_08DHFoOR;
R RWRH:RM0R#8F_Do
HOR
2;CRM8ObFlFMMC0
;
0C$bRVDC0CFPsR_0HN#Rs$sNRR5j0dFR2VRFR0HMCsoC;$
0bDCRCFV0P_Cs0R_.HN#Rs$sNRR5j04FR2VRFR0HMCsoC;k
VMHO0FbMRNH85R#:R0D8_FOoH_OPC0;FsR,I4RRI.:MRH0CCoss2RCs0kM0R#8F_Do_HOP0COFHsR#N
PsLHNDPCRN:sRR8#0_oDFHPO_CFO0s45I-84RF0IMF2Rj;C
Lo
HMRFRVsRR[HPMRNss'NCMoRFDFbR
RRVRHRR5[<I=R.02RERCM
RSRP5Ns[:2R=5RHHF'DI2+[;C
SD
#CSPRRN[s52=R:R''j;C
SMH8RVR;
R8CMRFDFbR;
R0sCkRsMP;Ns
8CMR8bN;k
VMHO0FoMRCI0_HE80_IU5HE80:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:R8IH0UE/;R
RH5VR58IH0lERFU8R2RR>c02RE
CMRRRRPRND:P=RN+DRR
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0I0H8E;_U
MVkOF0HMCRo0H_I8_0E.H5I8:0ER0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RDPNRR:=I0H8E;/.
sRRCs0kMNRPDC;
Mo8RCI0_HE80_
.;VOkM0MHFR0oC_8IH0IE5HE80RH:RMo0CCRs2skC0sDMRCFV0P_Cs0R_.HP#
NNsHLRDCPRND:CRDVP0FC0s__
.;LHCoMR
RP5ND4:2R=CRo0H_I8_0E.H5I820E;R
RH5VRI0H8EFRl8RR.=2RjRC0EMR
RRNRPD25jRR:=jR;
R#CDCR
RRNRPD25jRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCI0_HE80;k
VMHO0FoMRCI0_HE8058IH0:ERR0HMCsoC2CRs0MksRVDC0CFPsR_0HP#
NNsHLRDCPRND:CRDVP0FC0s_RR:=5Rj,jj,R,2Rj;C
Lo
HMRNRPD25dRR:=o_C0I0H8E5_UI0H8E
2;RNRO#5CRI0H8EFRl82RUR
H#RERICcMRRd|RRR=>P5ND.:2R=;R4
IRRERCM.>R=RDPN5R42:4=R;R
RIMECR=4R>NRPD25jRR:=4R;
RCIEM0RFE#CsRR=>MDkD;R
RCRM8OCN#;R
RskC0sPMRN
D;CRM8o_C0I0H8EO;
F0M#NRM0I0H8Es_NsRN$:CRDVP0FC0s_RR:=o_C0I0H8EH5I820E;F
OMN#0MI0RHE80_sNsNn$_cRR:D0CVFsPC_.0_RR:=o_C0I0H8EH5I820E;k
VMHO0FoMRCM0_k4l_.8U5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C04E/.
U;RVRHR855CEb0R8lFRU4.2RR>424.RC0EMR
RRNRPD=R:RDPNR4+R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._4UV;
k0MOHRFMo_C0D0CVFsPC_5nc80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF842.U;M
C8CRo0C_DVP0FCns_cV;
k0MOHRFMo_C0M_kln8c5CEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0RR<=4R4.NRM880CbERR>cRU20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kln
c;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_nV;
k0MOHRFMo_C0C_M880CbEH5#x:CRR0HMCsoCR8;RCEb0RH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDlCRH#M_HRxC:MRH0CCos=R:R
j;LHCoMR
Rl_HM#CHxRR:=80CbER;
RRHV5x#HCRR<80CbE02RE
CMRRRRl_HM#CHxRR:=#CHx;R
RCRM8H
V;RCRs0MksRMlH_x#HCC;
Mo8RCC0_M88_CEb0;-
-O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5855CEb0R4-R2RR/dR.2+5R55b8C0-ERRR42lRF8dR.2/nR42R2;R-R-RFyRVqR)vXd.4O1RC#DDRCMC8RC8
MOF#M0N0kRMlC_OD4D_.:URR0HMCsoCRR:=o_C0M_kl45.U80CbE
2;O#FM00NMRVDC0CFPsc_nRH:RMo0CC:sR=CRo0C_DVP0FCns_cC58b20E;F
OMN#0MM0RkOl_C_DDn:cRR0HMCsoCRR:=o_C0M_klnDc5CFV0P_Csn;c2
MOF#M0N0CRDVP0FCds_.RR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,ncR2nc;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bC4R.UHN#Rs$sNRk5MlC_OD4D_.8URF0IMF,RjR8IH04E-RI8FMR0FjF2RV0R#8F_Do;HO
b0$CkRF0k_L#$_0bnC_c#RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdH.R#sRNsRN$5lMk_DOCD._dRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO0;
$RbCF_k0L_k#0C$b_R4nHN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_k4#_.:URR0Fk_#Lk_b0$C._4UR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kn#_cRR:F_k0L_k#0C$b_;ncRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_Rd.:kRF0k_L#$_0bdC_.R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_k4#_nRR:F_k0L_k#0C$b_;4nRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C_DD4R.U8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDF_k0CnM_cRR:#_08DHFoO#;
HNoMDkRF0M_C_Rd.:0R#8F_Do;HO
o#HMRNDF_k0C4M_nRR:#_08DHFoO#;
HNoMDsRI0M_CR#:R0D8_FOoH_OPC05FsM_klODCD_U4.RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rnc:0R#8F_Do;HO
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F58nRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2F
OMN#0MD0R#IL_HE80RH:RMo0CC:sR=HRI8-0EUI*5HE80_sNsNd$522-4-Ic*HE80_sNsN.$52*-.I0H8Es_Ns5N$4I2-HE80_sNsNj$520;
$RbC0_lbNNss$HUR#sRNsRN$58IH0NE_s$sN5-d24FR8IFM0RRj2F#VR0D8_FOoH_OPC05Fs(FR8IFM0R;j2
o#HMRND0_lbU._d,lR0b__U4:nRRb0l_sNsN;$U
0N0skHL0\CR3lsN_VFV#\C0R#:R0MsHoL;
CMoH
R
RR-R-RRQVNs88I0H8ERR<(#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDI8_N8<sR=jR"jjjjj&"RR_N8s5Coj
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<"=Rjjjjj&"RR_N8s5Co4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjjj&"RR_N8s5Co.FR8IFM0R;j2
RRRR8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CRRRRRRRRD_FINs88RR<="jjj"RR&Ns8_Cdo5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
cSzSH:RVNR58I8sHE80R6=R2CRoMNCs0SC
SIDF_8N8s=R<Rj"j"RR&Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;z
S6RS:H5VRNs88I0H8ERR=no2RCsMCN
0CSFSDI8_N8<sR=jR''RR&Ns8_C6o5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRDRRFNI_8R8s<N=R8C_soR5n8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
n;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR(R:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rh7Q;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz
(;RRRRzRUR:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR=QR7hR;
RCRRMo8RCsMCNR0Cz
U;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRRg:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soR;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zg
RRRRjz4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C
o;RRRRCRM8oCCMsCN0Rjz4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR44RH:RVNR58_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,q)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRR8RN_osCRR<=q)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC4Rz4R;
RzRR4:.RRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);RRRRCRM8oCCMsCN0R.z4;R
RRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4RzdRR:VRFsHMRHRk5MlC_OD4D_.-URRR428MFI0jFRRMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:cRRRHV58N8s8IH0>ERRR(2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2R(RH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F(=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
c;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR46:VRHR85N8HsI8R0E<(=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRnz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vU4.RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloHC5*U4.2RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*U4.,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4R.U:)RXq.v4U1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRq6=D>RFNI_858s6R2,q=nR>FRDI8_N8ns52S,
SSSSSWRR >R=R0Is_5CMHR2,WiBpRR=>B,piR=mR>kRF0k_L#._4U,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k4#_.HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4RznR;
RRRRCRM8oCCMsCN0Rdz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0R4NRnFRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:(RRRHV5lMk_DOCDc_nR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4URH:RVNR58I8sHE80R(>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mc_nRR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;UN
RRRRRRRRUz4LRR:H5VRNs88I0H8ERR=(MRN8kRMlC_OD4D_.=URRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMn<cR=4R''ERIC5MR5_N8s5Con=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMn<cR= RWRCIEM5R5Ns8_Cno52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0RUz4LR;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:gRRRHV58N8s8IH0<ER=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rnc<'=R4
';RRRRRRRRRRRRRRRRI_s0CnM_c=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RzgR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
SRzRRO_E	.RR:H5VRI0H8Es_Ns_N$n4c52RR>jo2RCsMCN
0CRRRRRRRRzR.j:FRVsRR[H5MRI0H8Es_Ns_N$n4c52RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERR[.*R.-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*;[2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:Xv)qn.cX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R74=H>RMC_soH5I8-0E.-*[4R2,7=jR>MRH_osC58IH0.E-*.[-2q,Rj>R=RIDF_8N8s25j,4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FINs885,d2RRqc=D>RFNI_858scR2,q=6R>FRDI8_N86s52S,
SSSSSWRR >R=R0Is__CMnRc,WiBpRR=>B,piRRm4=F>RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.-*[4R2,m=jR>kRF0k_L#c_n5lMk_DOCDc_n,8IH0.E-*.[-2
2;RRRRRRRRRRRRRRRRF_k0s5CoI0H8E*-.[2-4RR<=F_k0L_k#nMc5kOl_C_DDnIc,HE80-[.*-R42IMECRk5F0M_C_Rnc=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC58IH0.E-*.[-2=R<R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.[2-.RCIEMFR5kC0_Mc_nR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.j
RSSCRM8oCCMsCN0REzO	;_.
RSSz	OE_:4RRRHV58IH0NE_s$sN_5ncj>2RRRj2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4U&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRI.*HE80_sNsNn$_c254R4-R2RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URR,ncRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80R.-R*8IH0NE_s$sN_5nc4;22
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)nqvcRR:)nqvc1X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5CoI0H8E*-.I0H8Es_Ns_N$n4c522-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52q,R6>R=RIDF_8N8s256,S
SSSSSR RWRR=>I_s0CnM_cW,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5ncM_klODCD_,ncI0H8E*-.I0H8Es_Ns_N$n4c522-42R;
RRRRRRRRRRRRRFRRks0_CIo5HE80-I.*HE80_sNsNn$_c254-R42<F=RkL0_kn#_ck5MlC_ODnD_cH,I8-0E.H*I8_0ENNss$c_n5-424I2RERCM50Fk__CMn=cRR''42DRC#'CRZ
';RRRRRRRRR8CMRMoCC0sNCORzE4	_;R
RRSRRR8CMRMoCC0sNC4Rz(R;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR.4:VRHRk5MlC_ODdD_.RR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.z.NRR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''42MRN8NR58C_so256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN..;R
RRRRRR.Rz.:LRRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn/cR=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=RjR'2NRM85_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rz.
L;RRRRRRRRzO..RH:RVNR58I8sHE80R(=RR8NMRlMk_DOCDc_nR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRN558C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5Ns8_Cno52RR='24'R8NMR85N_osC5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.O
RRRRRRRR.z.8RR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODnD_c=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI06FR2RR=M_klODCD_2nc2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR62=kRMlC_ODnD_cR22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;.8
RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.d
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CSRRRREzO	R_U:VRHRH5I8_0ENNss$25dRj>R2CRoMNCs0SC
SEzO	C_D6RR:H5VRI0H8E=R>RIU*HE80_sNsNd$52MRN8HRI8R0E>U=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8M5H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_.25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0R8IH0DE-#IL_HE80RMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdH.,[<2R=lR0b__Udj.52[5H-8IH0DE+#IL_HE802R;
RRRRRRRRRRRRRRRRR0Fk_osC52H[RR<=F_k0L_k#dM.5kOl_C_DDdH.,[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';SSSSCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRRUz.RV:RF[sRRRHMI0H8Es_Ns5N$d42-RI8FMR0F4CRoMNCs0RC
RRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNCH5I8R0E-#RDLH_I8R0E-*R[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0-ERR-5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vRd.:)RXq.vdXRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_CIo5HE80-LD#_8IH0UE-*([+RI8FMR0FI0H8E#-DLH_I8-0EU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SRSSRNRR#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#dM.5kOl_C_DDdI.,HE80-LD#_8IH0UE-*H[+[<2R=lR0b__Ud[.52[5H2R;
RRRRRRRRRRRRRRRRR0Fk_osC58IH0DE-#IL_HE80-[U*+2H[RR<=F_k0L_k#dM.5kOl_C_DDdI.,HE80-LD#_8IH0UE-*H[+[I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzED	_C
6;SOSzEo	_0:6RRRHV58IH0>ER=RRUNRM8I0H8EFRl8RRU>6=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8E&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vRd.:)RXq.vdX
U1SRSSRbRRFRs0lRNb5=7R>NRb8M5H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_dU_.H5I8_0ENNss$25d-242;S
SS#SN#MHoRV:RFHsR[MRHR8IH04E-RI8FMR0FI0H8E#-DLH_I8R0EoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.H5I8_0ENNss$25d-542HI[-HE80+LD#_8IH0;E2
RRRRRRRRRRRRRRRRFRRks0_CHo5[<2R=kRF0k_L#._d5lMk_DOCD._d,2H[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMR;
RRRRRRRRRzRR.:URRsVFRH[RMHRI8_0ENNss$25d-8.RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC*5[U&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5+5[4U2*2R;
RRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRqz)vRd.:)RXq.vdXRU1
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_CUo5*([+RI8FMR0FU2*[,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piR=mR>lR0b__Ud[.52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_5d.M_klODCD_,d.U+*[HR[2<0=RlUb__5d.[H25[
2;RRRRRRRRRRRRRRRRRkRF0C_so*5U[[+H2=R<R0Fk_#Lk_5d.M_klODCD_,d.U+*[HR[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	o;06
zSSO_E	MRR:H5VRI0H8ERR<Uo2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC25U;R
RRRRRRRRRRCRLo
HMSRSRR)Rzq.vdRX:R)dqv.1XU
SSSRRRRb0FsRblNRR57=b>RNH85MC_soH5I8-0E4FR8IFM0R8IH0DE-#IL_HE802U,R,#RDLH_I8-0E4R2,q=jR>FRDI8_N8js52S,
SSSSSqRR4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2RRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__Udj.52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFRRjoCCMsCN0
SSSSFRRkL0_kd#_.k5MlC_ODdD_.[,H2=R<Rb0l_dU_.25j52H[;R
RRRRRRRRRRRRRRRRRF_k0s5CoHR[2<F=RkL0_kd#_.k5MlC_ODdD_.[,H2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''S;
SCSSMo8RCsMCNR0CNH##o
M;SMSC8CRoMNCs0zCRO_E	MS;
S8CMRMoCC0sNCORzEU	_;S
Sz	OE_:cRRRHV58IH0NE_s$sN5R.2>2RjRMoCC0sNCR
RRRRRR.RzcR_c:VRHRH5I8R0E>c=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=H>RMC_so25d,.R7RR=>HsM_C.o527,R4>R=R_HMs5Co4R2,7=jR>MRH_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,q=cR>FRDI8_N8cs52W,R >R=R0Is__CMdR.,WiBpRR=>B,piRS
SSSSSRdRmRR=>F_k0L_k#dM.5kOl_C_DDdd.,2m,R.>R=R0Fk_#Lk_5d.M_klODCD_,d..
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,,42RRmj=F>RkL0_kd#_.k5MlC_ODdD_.2,j2R;
RRRRRRRRRRRRRFRRks0_Cdo52=R<R0Fk_#Lk_5d.M_klODCD_,d.dI2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5R42<F=RkL0_kd#_.k5MlC_ODdD_.2,4RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.ccR;
RRRRRzRR.dc_RH:RVIR5HE80Rd=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq.vdRD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*n2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo5;c2
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR)dqv.RR:Xv)qdc.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d='>RjR',7=.R>MRH_osC5,.2RR74=H>RMC_so254,jR7RR=>HsM_Cjo52S,
SRSRRRRRRRRRRRRRq=jR>FRDI8_N8js52q,R4>R=RIDF_8N8s254,.RqRR=>D_FINs885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8N8s25d,cRqRR=>D_FINs885,c2RRW =I>RsC0_M._d,BRWp=iR>pRBi
,RSSSSSRSRm=dR>bRFCRM,m=.R>kRF0k_L#._d5lMk_DOCD._d,,.2
SSSSRSSRRm4=F>RkL0_kd#_.k5MlC_ODdD_.2,4,jRmRR=>F_k0L_k#dM.5kOl_C_DDdj.,2
2;RRRRRRRRRRRRRRRRF_k0s5Co.<2R=kRF0k_L#._d5lMk_DOCD._d,R.2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5R42<F=RkL0_kd#_.k5MlC_ODdD_.2,4RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so25jRR<=F_k0L_k#dM.5kOl_C_DDdj.,2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz_.cdS;
S8CMRMoCC0sNCORzEc	_;S
Sz	OE_:.RRRHV58IH0NE_s$sN5R42>2RjRMoCC0sNCR
RRRRRR.RzcRR:VRFs[MRHRH5I8_0ENNss$254R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*8IH0NE_s$sN5-d2.-*[.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0UE-*8IH0NE_s$sN5-d2.2*[;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRv)qd..X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7j=H>RMC_soH5I8-0EUH*I8_0ENNss$25d-[.*-,.2RR74=H>RMC_soH5I8-0EUH*I8_0ENNss$25d-[.*-,42RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m=jR>kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*8IH0NE_s$sN5-d2.-*[.
2,SSSSSRSRm=4R>kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*8IH0NE_s$sN5-d2.-*[4;22
RRRRRRRRRRRRRRRR0Fk_osC58IH0UE-*8IH0NE_s$sN5-d2.-*[4<2R=kRF0k_L#._d5lMk_DOCD._d,8IH0UE-*8IH0NE_s$sN5-d2.-*[4I2RERCM50Fk__CMd=.RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5CoI0H8E*-UI0H8Es_Ns5N$d.2-*.[-2=R<R0Fk_#Lk_5d.M_klODCD_,d.I0H8E*-UI0H8Es_Ns5N$d.2-*.[-2ERIC5MRF_k0CdM_.RR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.c
CSSMo8RCsMCNR0Cz	OE_
.;SOSzE4	_RH:RVIR5HE80_sNsNj$52RR>jo2RCsMCN
0CRRRRRRRRzR.c:VRHRH5I8R0ElRF8URR=4o2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*c&2RR""WRH&RMo0CCHs'lCNo5Rj2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+dR.,80CbER22&XR""RR&HCM0o'CsHolNC254;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRv)qd4.X1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52q,Rc>R=RIDF_8N8s25c, RWRR=>I_s0CdM_.W,RBRpi=B>RpRi,m>R=R0Fk_#Lk_5d.M_klODCD_,d.j;22
RRRRRRRRRRRRRRRR0Fk_osC5Rj2<F=RkL0_kd#_.k5MlC_ODdD_.2,jRCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.
c;SMSC8CRoMNCs0zCRO_E	4R;
RCRRMo8RCsMCNR0Cz;.4RRRRRRRRR
R
RRRR-t-RCsMCNR0CNnR4RsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR.Rz6RR:H5VRM_klODCD_R4n=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR62M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR.RnN:VRHR85N8HsI8R0E>RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='24'R8NMR85N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''42MRN8NR58C_so256R'=R4R'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzn
N;RRRRRRRRzL.nRH:RVNR58I8sHE80R(>RR8NMRlMk_DOCDc_nR4=RR8NMRlMk_DOCD._dRj=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RR(2=kRMlC_OD4D_.RU2NRM85_N8s5Con=2RR''42MRN8NR58C_so256R'=RjR'2NRM85_N8s5Coc=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='2j'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nL
RRRRRRRRnz.ORR:H5VRNs88I0H8ERR>(MRN8kRMlC_ODnD_cRR=jMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_CNo58I8sHE80-84RF0IMF2R(RM=RkOl_C_DD42.UR8NMR85N_osC5Rn2=jR''N2RM58RNs8_C6o52RR='24'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=RjR'2NRM85_N8s5Co6=2RR''42MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO.n;R
RRRRRR.Rzn:8RRRHV58N8s8IH0>ERRN(RMM8RkOl_C_DDn=cRRNjRMM8RkOl_C_DDd=.RRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0(FR2RR=M_klODCD_U4.2MRN8NR58C_so25nR'=RjR'2NRM85_N8s5Co6=2RR''j2MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC58N8s8IH04E-RI8FMR0F(=2RRlMk_DOCD._4UN2RM58RNs8_Cno52RR='2j'R8NMR85N_osC5R62=jR''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.8R;
RRRRRzRR.RnC:VRHR85N8HsI8R0E=RR(NRM8M_klODCD_Rnc=RR4NRM8M_klODCD_Rd.=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM585N_osC5Rn2=4R''N2RM58RNs8_C6o52RR='24'R8NMR85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5Con=2RR''42MRN8NR58C_so256R'=R4R'2NRM8R85N_osC5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;nC
RRRRRRRRnz.VRR:H5VRNs88I0H8ERR=(MRN8kRMlC_ODnD_cRR=4MRN8kRMlC_ODdD_.RR=jo2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5Ns8_Cno52RR='24'R8NMR85N_osC5R62=jR''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRN558C_so25nR'=R4R'2NRM85_N8s5Co6=2RR''j2MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzV.n;R
RRRRRR.Rzn:oRRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn=cRRNjRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR5_N8s5Co6=2RR''42MRN8NR58C_so25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM585N_osC5R62=4R''N2RM58RNs8_Cco52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.oR;
RRRRRzRR.RnE:VRHR85N8HsI8R0E=RR6NRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRN558C_so85N8HsI8-0E4FR8IFM0RRc2=kRMlC_ODdD_.R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR5_N8s5CoNs88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rnz.ER;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:(RRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.Rz(R;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
SRzRRO_E	URR:H5VRI0H8Es_Ns5N$d>2RRRj2oCCMsCN0
zSSO_E	DRC6:VRHRH5I8R0E>U=R*8IH0NE_s$sN5Rd2NRM8I0H8E=R>RRU2oCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)q4:nRRLDNCHDR#1R"1Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*2d.R"&RW&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE802RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0+ERR;U2
RRRRRRRRRRRRoLCHSM
SRRRRqz)vR4n:)RXqnv4X
U1SRSSRbRRFRs0lRNb5=7R>NRb8M5H_osC58IH04E-RI8FMR0FI0H8E#-DLH_I820E,,RURLD#_8IH04E-2q,Rj>R=RIDF_8N8s25j,S
SSSSSR4RqRR=>D_FINs885,42RRq.=D>RFNI_858s.R2,q=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,pi
SSSSRSSR=mR>lR0b__U4jn52
2;SSSSNH##o:MRRsVFRRH[HIMRHE80-84RF0IMFHRI8-0ED_#LI0H8ECRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nHR[2<0=RlUb__54njH25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRRkRF0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHR8IH0NE_s$sN5-d24FR8IFM0Ro4RCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCI0H8ERR-D_#LI0H8ERR-54[-22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)q4:nRRqX)vX4nU
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_soH5I8-0ED_#LI0H8E*-U[R+(8MFI0IFRHE80-LD#_8IH0UE-*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>lR0b__U4[n52
2;SRSSRNRR#o#HMRR:VRFsHH[RMRR(8MFI0jFRRMoCC0sNCS
SSRSRF_k0L_k#4Mn5kOl_C_DD4In,HE80-LD#_8IH0UE-*H[+[<2R=lR0b__U4[n52[5H2R;
RRRRRRRRRRRRRRRRR0Fk_osC58IH0DE-#IL_HE80-[U*+2H[RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-LD#_8IH0UE-*H[+[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRCRM8oCCMsCN0R#N#H;oM
RRRRRRRRRRRR8CMRMoCC0sNC.RzUS;
S8CMRMoCC0sNCORzED	_C
6;SOSzEo	_0:6RRRHV58IH0>ER=RRUNRM8I0H8EFRl8RRU>6=R2CRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0-ERRLD#_8IH0RE2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.d+.RR,4nRb8C02E2R"&RX&"RR0HMCsoC'NHloIC5HE80RD-R#IL_HE80RU+R2R;
RRRRRRRRRLRRCMoH
RSSRzRR)4qvnRR:Xv)q4UnX1S
SSRRRRsbF0NRlb7R5RR=>b5N8HsM_CIo5HE80-84RF0IMFHRI8-0ED_#LI0H8ER2,UD,R#IL_HE80-,42RRqj=D>RFNI_858sj
2,SSSSSRSRq=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,dRqRR=>D_FINs885,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBiS,
SSSSSmRRRR=>0_lbUn_458IH0NE_s$sN5-d24;22
SSSS#N#HRoM:FRVs[RHRRHMI0H8ER-48MFI0IFRHE80-LD#_8IH0oERCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_458IH0NE_s$sN5-d24H25[H-I8+0ED_#LI0H8E
2;RRRRRRRRRRRRRRRRRkRF0C_so[5H2=R<R0Fk_#Lk_54nM_klODCD_,4nHR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
SSSS8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRR.RzURR:VRFs[MRHR8IH0NE_s$sN5-d2.FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oC[2*UR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC54[+22*U;R
RRRRRRRRRRRRRLHCoMR
RRRRRRRRRRRRRzv)q4:nRRqX)vX4nU
1RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so*5U[R+(8MFI0UFR*,[2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>lR0b__U4[n52
2;SSSSNH##o:MRRsVFRRH[H(MRRI8FMR0FjCRoMNCs0SC
SRSSR0Fk_#Lk_54nM_klODCD_,4nU+*[HR[2<0=RlUb__54n[H25[
2;RRRRRRRRRRRRRRRRRkRF0C_so*5U[[+H2=R<R0Fk_#Lk_54nM_klODCD_,4nU+*[HR[2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR8CMRMoCC0sNC#RN#MHo;R
RRRRRRRRRRMRC8CRoMNCs0zCR.
U;SMSC8CRoMNCs0zCRO_E	o;06
zSSO_E	MRR:H5VRI0H8ERR<Uo2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCU
2;RRRRRRRRRRRRLHCoMS
SRRRRzv)q4:nRRqX)vX4nUS1
SRSRRFRbsl0RN5bR7>R=R8bN5_HMs5CoI0H8ER-48MFI0IFRHE80-LD#_8IH0,E2RRU,D_#LI0H8E2-4,jRqRR=>D_FINs885,j2
SSSSRSSRRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52q,Rd>R=RIDF_8N8s25d, RWRR=>I_s0C4M_nW,RBRpi=B>Rp
i,SSSSSRSRm>R=Rb0l_4U_n25j2S;
SNSS#o#HMRR:VRFsHH[RMHRI8-0E4FR8IFM0RojRCsMCN
0CSSSSRkRF0k_L#n_45lMk_DOCDn_4,2H[RR<=0_lbUn_455j2H;[2
RRRRRRRRRRRRRRRRFRRks0_CHo5[<2R=kRF0k_L#n_45lMk_DOCDn_4,2H[RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;S
SSMSC8CRoMNCs0NCR#o#HMS;
S8CMRMoCC0sNCORzEM	_;S
SCRM8oCCMsCN0REzO	;_U
zSSO_E	cRR:H5VRI0H8Es_Ns5N$.>2RRRj2oCCMsCN0
RRRRRRRRgz._:cRRRHV58IH0>ER=2RcRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC25c;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q4cnX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5R7d=H>RMC_so25d,.R7RR=>HsM_C.o527,R4>R=R_HMs5Co4R2,7=jR>MRH_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,SR
SSSSSmRRd>R=R0Fk_#Lk_54nM_klODCD_,4ndR2,m=.R>kRF0k_L#n_45lMk_DOCDn_4,,.2
SSSSRSSRRm4=F>RkL0_k4#_nk5MlC_OD4D_n2,4,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4jn,2
2;RRRRRRRRRRRRRRRRF_k0s5Cod<2R=kRF0k_L#n_45lMk_DOCDn_4,Rd2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5R.2<F=RkL0_k4#_nk5MlC_OD4D_n2,.RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so254RR<=F_k0L_k#4Mn5kOl_C_DD44n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cjo52=R<R0Fk_#Lk_54nM_klODCD_,4njI2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0Rgz._
c;RRRRRRRRz_.gdRR:H5VRI0H8ERR=do2RCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)4qvnRR:DCNLD#RHR1"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_U4.*U4.RM+RkOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25jR"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCD._4U.*4URR+M_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oCc
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)Rzqnv4R):Rqnv4XRc1
RRRRRRRRRRRRRRRRsbF0NRlb7R5d>R=R''j,.R7RR=>HsM_C.o527,R4>R=R_HMs5Co4R2,7=jR>MRH_osC5,j2
SSSRRRRRRRRRRRRRjRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,SR
SSSSSmRRd>R=RCFbMm,R.>R=R0Fk_#Lk_54nM_klODCD_,4n.
2,SSSSSRSRm=4R>kRF0k_L#n_45lMk_DOCDn_4,,42RRmj=F>RkL0_k4#_nk5MlC_OD4D_n2,j2R;
RRRRRRRRRRRRRFRRks0_C.o52=R<R0Fk_#Lk_54nM_klODCD_,4n.I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4<2R=kRF0k_L#n_45lMk_DOCDn_4,R42IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5Rj2<F=RkL0_k4#_nk5MlC_OD4D_n2,jRCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRMRC8CRoMNCs0zCR.dg_;S
SCRM8oCCMsCN0REzO	;_c
zSSO_E	.RR:H5VRI0H8Es_Ns5N$4>2RRRj2oCCMsCN0
RRRRRRRRjzdRV:RF[sRRRHM58IH0NE_s$sN5R42-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a11"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo58IH0UE-*8IH0NE_s$sN5-d2.-*[.&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNCH5I8-0EUH*I8_0ENNss$25d-[.*2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n.
1RRRRRRRRRRRRRRRRRb0FsRblNRj57RR=>HsM_CIo5HE80-IU*HE80_sNsNd$52*-.[2-.,4R7RR=>HsM_CIo5HE80-IU*HE80_sNsNd$52*-.[2-4,jRqRR=>D_FINs885,j2RRq4=D>RFNI_858s4R2,q=.R>FRDI8_N8.s52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFNI_858sdR2,W= R>sRI0M_C_,4nRpWBi>R=RiBp,jRmRR=>F_k0L_k#4Mn5kOl_C_DD4In,HE80-IU*HE80_sNsNd$52*-.[2-.,S
SSSSSR4RmRR=>F_k0L_k#4Mn5kOl_C_DD4In,HE80-IU*HE80_sNsNd$52*-.[2-42R;
RRRRRRRRRRRRRFRRks0_CIo5HE80-IU*HE80_sNsNd$52*-.[2-4RR<=F_k0L_k#4Mn5kOl_C_DD4In,HE80-IU*HE80_sNsNd$52*-.[2-4RCIEMFR5kC0_Mn_4R'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soH5I8-0EUH*I8_0ENNss$25d-[.*-R.2<F=RkL0_k4#_nk5MlC_OD4D_nH,I8-0EUH*I8_0ENNss$25d-[.*-R.2IMECRk5F0M_C_R4n=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNCdRzjS;
S8CMRMoCC0sNCORzE.	_;S
Sz	OE_:4RRRHV58IH0NE_s$sN5Rj2>2RjRMoCC0sNCR
RRRRRRdRz4RR:H5VRI0H8EFRl8RRU=2R4RMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"1aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_OD4D_.4U*.+URRlMk_DOCDc_n*Rnc+kRMlC_ODdD_..*d2RR&"RW"&MRH0CCosl'HN5oCj&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C0ME5kOl_C_DD4*.U4R.U+kRMlC_ODnD_cc*nRM+RkOl_C_DDdd.*.RR+4Rn,80CbER22&XR""RR&HCM0o'CsHolNC254;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q44nX1RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,j2RRqj=D>RFNI_858sjR2,q=4R>FRDI8_N84s52q,R.>R=RIDF_8N8s25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDI8_N8ds52W,R >R=R0Is__CM4Rn,WiBpRR=>B,piR=mR>kRF0k_L#n_45lMk_DOCDn_4,2j2;R
RRRRRRRRRRRRRRkRF0C_so25jRR<=F_k0L_k#4Mn5kOl_C_DD4jn,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;d4
CSSMo8RCsMCNR0Cz	OE_
4;RRRRR8CMRMoCC0sNC.Rz6R;RRRRRRRRR
M
C8sRNO0EHCkO0s#CRCODC0N_sl
;

