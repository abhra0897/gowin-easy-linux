-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRR:wRRH8GC-HbFMb0RNNO	o5CRtCCMsRHOb	NONRoC8DCON0sNH2FM
R--RRRRRRRRRRRR:-
-RpRRHNLssR$RRR:Ra#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRRR:R#L$lFODHN$DDRlMNCQ8R 3  
R--RRRRRRRRRRRR:-
-R7RRCDPCFsbC#R:RqCOODsDCN]Re7ap-BMRN8 RQ u R4nj(RsWF	oHMRFtsk-b
-RRRRRRRRRRRR
R:-R-RRsukbCF#R:RRRERaHb#RNNO	oRC#8HCVMRC#LHN#OHRLM$NsRGVHCb8RF0HM
R--RRRRRRRRRRRR:NRRsEH0lHC0OkRVMHO0F
M#-R-RRRRRRRRRR:RR
R--RFRh0RCRRRRR:aRRERH#b	NONRoClRN$LlCRFV8HHRC80HFRMkOD8NCR808HHNFMDNR80-N
-RRRRRRRRRRRRRR:RJsCkCHs8$RLRF0FDR#,LRk0Hl0RkR#0HMMRFNRI$ERONCMoRC0E
R--RRRRRRRRRRRR:CRRGs0CMRNDHCM0sOVNCF#RsHR#lNkD0MHFRELCNFPHsVRFRC0E
R--RRRRRRRRRRRR:8RRCs#OHHb0FRM3QH0R#CRbs#lH#DHLCFR0R8N8RlOFl0CM#MRN8s/F
R--RRRRRRRRRRRR:NRR0H0sLCk0#FR0RC0ERObN	CNoRO8CDNNs0MHF#L,RkM0RF00RFERONCMo
R--RRRRRRRRRRRR:FRRsCR8DCC0R$NMRHFsoNHMDHRDMRC#F0VREbCRNNO	o8CRCNODsHN0F
M3-R-RRRRRRRRRR:RRRERaCNRbOo	NCFRL8l$RNL$RCERONCMo8MRFDH$RMORNO8FsNCMOR0IHE-
-RRRRRRRRRRRRRR:R0REC0lCs#VRFRNBDkR#C4FnRVER0H##R08NMN3s8
R--RRRRRRRRRRRR:-
-R---------------------------------------------------------------------
-RCf)PHH#FRM:4j..R-f
-7RfN:0CRj.jUc-j-R4j44(:ng:jRg+jd5jRa,EkRR4jqRbs.Ujj2
Rf---R-----------------------------------------------------------------
--
Ck#R71a3Xa a3QmN;DD
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   3vhz B)Q_71a3DND;#
kC RQ V 3H8GC_FVDN00_$#bC3DND;b

NNO	oVCRH8GC_MoCCOsH_ob	R
H#RCRoMHCsO
R5RRRR-)-RF8kMHRMos0FkHRMC0kFR#HCRMHRVGRC8bMFH0V,RH8GC_ksFMF8RsHRVG_C80MskOCN0
RRRRGVHCs8_F8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM;R
RR-R-RCmPsFVDIFRskM0HCFR0RCk#RRHMVCHG8FRbH,M0RGVHC#8_Ns0kNR0CFVsRH8GC_NIsbR
RRHRVG_C8FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8#kN0sCN0;R
RR-R-R0 GsLNRHR0#k8#CRRHM8HHP8sCRFHk0M
C#RRRRVCHG8k_oN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=dR;
R-RR-VRQRza) 0,RERCM0MksRVFVRsINMoHM#MRFR""XRFbsbNNo0MHF
RRRR_MFIMNsHRMoRRRRRRRRRRR:Apmm RqhRRRRRRRRRRRRRRRRR=R:RDVN#RC
R2RR;R

RR--qEk0F7sRN8PHR#AHERFb5H8L#bEF@E@P8FD3s
o2RFROMN#0MB0RF)b$H0oEhHF0O:CRR)1aQRht:R=
R"RRB$FbsEHo0jR.jLUR$ RQ R 3qRDDsEHo0s#RCs#CP3C8"
;
R-R-R#LNCMRz#MHoCV8RH8GCRHbFM00R$,bCRI8FMR0F8CHsOF0HM#RN#Ckl8R
R0C$bR)zh p1me_ 7kGVHCH8R#sRNsRN$5aQh )t RMsNo<CR>F2RVaR17p_zmBtQ;R
R-L-RNR#C1MHoCV8RH8GCRHbFM00R$,bCRI8FMR0F8CHsOF0HM#RN#Ckl8R
R0C$bR)zh p1me_ 7#GVHCH8R#sRNsRN$5aQh )t RMsNo<CR>F2RVaR17p_zmBtQ;R

RHNDNz#R_HkVGRC8Hz#Rh1) m pe7V_kH8GC;R
RNNDH#_Rz#GVHCH8R#hRz)m 1p7e _H#VG;C8
R
R#0kL$RbCkGVHCH8R#CRs#PFDCz8Rh1) m pe7V_kH8GC;R
R#0kL$RbC#GVHCH8R#CRs#PFDCz8Rh1) m pe7V_#H8GC;R

R=--=========================================================================R=
RR--q0sHE0lCHmORbNCs0#Fs:R
R-=-==========================================================================R

RR--qFL#DCk0RDPNkRC,.R'#ObFlDCClMR0
RR--NRL##GVHCN85RI8FMR0FL=2RRH#VG5C8NR+48MFI0LFR2R
RVOkM0MHFRL"N#5"RNRso:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RohCNF0HM.,R'O#RFDlbCMlC0R
R---RRH#VG5C8NFR8IFM0RRL2=VR#H8GC54N+RI8FMR0FLR2
RMVkOF0HM-R""NR5s:oRR)zh p1me_ 7#GVHCs82Cs0kMhRz)m 1p7e _H#VG;C8
R
R-q-R808HH
FMR-R-RHkVG5C8NFR8IFM0RRL2+VRkH8GC58ORF0IMF2R8
-RR-RRR=VRkH8GC5GlNHllk5ON,2R+48MFI0lFRHlMHkLl5,282
VRRk0MOHRFM"R+"5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-#-RVCHG8R5N8MFI0LFR2RR+#GVHCO85RI8FMR0F8R2
RR--RRR=#GVHCl85NlGHkNl5,+O24FR8IFM0RMlHHllk58L,2R2
RMVkOF0HM+R""DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RL1k0OsN0MHF
-RR-VRkH8GC58NRF0IMF2RLRk-RVCHG8R5O8MFI08FR2R
R-R-RRk=RVCHG8N5lGkHll,5NO42+RI8FMR0FlHHMl5klL2,82R
RVOkM0MHFR""-R,5DR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--#GVHCN85RI8FMR0FL-2RRH#VG5C8OFR8IFM0R
82R-R-R=RRRH#VG5C8lHNGl5klN2,O+84RF0IMFHRlMkHll,5L8
22RkRVMHO0F"MR-5"RDs,RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHC
8;
-RR-kRvDb0HDNHO0MHF
-RR-VRkH8GC58NRF0IMF2RLRk*RVCHG8R5O8MFI08FR2RR=kGVHCN85+4O+RI8FMR0FL2+8
VRRk0MOHRFM"R*"5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-#-RVCHG8R5N8MFI0LFR2RR*#GVHCO85RI8FMR0F8=2RRH#VG5C8N++O4FR8IFM0R8L+2R
RVOkM0MHFR""*R,5DR:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

RR--7HHP#MHF
-RR-VRkH8GC58NRF0IMF2RLRk/RVCHG8R5O8MFI08FR2RR=kGVHCN85-88RF0IMF-RLO2-4
VRRk0MOHRFM"R/"5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-#-RVCHG8R5N8MFI0LFR2RR/#GVHCO85RI8FMR0F8=2RRH#VG5C8N+-84FR8IFM0ROL-2R
RVOkM0MHFR""/R,5DR:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

RR--)NClHCM8sR
R-k-RVCHG8NR5RI8FMR0FLs2RCklRVCHG8OR5RI8FMR0F8R2
RR--RRR=kGVHC58RlHHMl5klN2,ORI8FMR0FlHHMl5klL2,82R
RVOkM0MHFRC"sl5"RDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VR#H8GCRR5N8MFI0LFR2CRslVR#H8GCRR5O8MFI08FR2R
R-R-RR#=RVCHG8lR5HlMHkNl5,RO28MFI0lFRHlMHkLl5,282
VRRk0MOHRFM"lsC"DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-R8vFk
DFR-R-RHkVGRC858NRF0IMF2RLR8lFRHkVGRC858ORF0IMF2R8
-RR-RRRRRRRRk=RVCHG8lR5HlMHkNl5,RO28MFI0lFRHlMHkLl5,2R82R
RVOkM0MHFRF"l85"RDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VR#H8GCRR5N8MFI0LFR2FRl8VR#H8GCRR5O8MFI08FR2R
R-R-RRRRRRRR=#GVHC58ROFR8IFM0RMlHHllk5RL,8
22RkRVMHO0F"MRl"F8R,5DR:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

R----------------------------------------------------------------------------R
R-Q-RMER0CR#Cs0FkH#MCRC0ERC"sNRD"F"sRMkN0s"NDRM5H0CCosR2
RR--NRsCOPFMCCs08MRH0NFRRGVHCb8RF0HMRlMkLRCsNRM80MECRC0ERCFbsHN0FHMR#R
R-b-RCFsVs8lC3QRR0#RHR#N#k8lCRN0E0ER0CsRNsRN$IDHDRRLCDoNsCMRCFEko3R
R-Q-RVER0CMRHbRk0H"#RsDCN"ER0C0MREsCRCRNDMLklCHsR#FROMsPC0RC8HFM0RVNRH8GCR
FVR-R-RC0ERl#NCHR#xNCR#ER0CHRVGRC8bMFH0MRHb3k0RVRQRC0ERlMkLRCsHN#RMHR"Mo0CC
s"R-R-RC0EM0RHRRH#OPFMCCs08MRH0VFRH8GCR0IHEER0CNRsMRoC5ED'HRoE8MFI0jFR2R3
R----------------------------------------------------------------------------R

RR--kGVHCN85RI8FMR0FL+2RRHkVG5C8NFR8IFM0RRL2=VRkH8GC54N+RI8FMR0FLR2
RMVkOF0HM+R""DR5Rz:Rh1) m pe7V_kH8GC;RRs: R)qRp2skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCO85RI8FMR0F8+2RRHkVG5C8OFR8IFM0RR82=VRkH8GC54O+RI8FMR0F8R2
RMVkOF0HM+R""DR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCN85RI8FMR0FL+2RRHkVG5C8NFR8IFM0RRj2=VRkH8GC54N+RI8FMR0FlHHMl5klj2,L2R
RVOkM0MHFR""+RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58NRF0IMF2RjRk+RVCHG8R5O8MFI08FR2RR=kGVHCO85+84RF0IMFHRlMkHll,5j8
22RkRVMHO0F"MR+5"RDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCN85RI8FMR0FL-2RRHkVG5C8NFR8IFM0RRL2=VRkH8GC54N+RI8FMR0FLR2
RMVkOF0HM-R""DR5Rz:Rh1) m pe7V_kH8GC;RRs: R)qRp2skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCO85RI8FMR0F8-2RRHkVG5C8OFR8IFM0RR82=VRkH8GC54O+RI8FMR0F8R2
RMVkOF0HM-R""DR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCN85RI8FMR0FL-2RRHkVG5C8NFR8IFM0RRj2=VRkH8GC54N+RI8FMR0FlHHMl5klj2,L2R
RVOkM0MHFR""-RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58NRF0IMF2RjRk+RVCHG8R5O8MFI08FR2RR=kGVHCO85+84RF0IMFHRlMkHll,5j8
22RkRVMHO0F"MR-5"RDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHCN85RI8FMR0FL*2RRHkVG5C8NFR8IFM0RRL2=VRkH8GC5+.N4FR8IFM0R2.L
VRRk0MOHRFM"R*"5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58ORF0IMF2R8Rk*RVCHG8R5O8MFI08FR2RR=kGVHC.85OR+48MFI0.FR8R2
RMVkOF0HM*R""DR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R

RR--kGVHC58RNFR8IFM0RRL2*VRkH8GCRR5N8MFI0jFR2RR=kGVHC58R.4N+RI8FMR0FLR2
RMVkOF0HM*R""DR5Rz:Rh1) m pe7V_kH8GC;RRs:qRhaqz)ps2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-k-RVCHG8NR5RI8FMR0FL*2RRHkVGRC858NRF0IMF2RjRk=RVCHG8.R5NR+48MFI0LFR2R
RVOkM0MHFR""*RR5D:qRhaqz)ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58NRF0IMF2RLRk/RVCHG8R5N8MFI0LFR2RR=kGVHCN85-8LRF0IMF-RLN2-4
VRRk0MOHRFM"R/"5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58NRF0IMF2RLRk/RVCHG8R5N8MFI0LFR2RR=kGVHCN85-8LRF0IMF-RLN2-4
VRRk0MOHRFM"R/"5:DRRq) ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GC58NRF0IMF2RLRk/RVCHG8R5N8MFI0jFR2RR=kGVHCN85RI8FMR0FL--N4R2
RMVkOF0HM/R""DR5Rz:Rh1) m pe7V_kH8GC;RRs:qRhaqz)ps2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-k-RVCHG8R5O8MFI0jFR2RR/kGVHCO85RI8FMR0F8=2RRHkVG5C8OR-88MFI0-FRO2-4
VRRk0MOHRFM"R/"5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8
;
R-R-RHkVGRC858NRF0IMF2RLRlsCRHkVGRC858NRF0IMF2RLRk=RVCHG8NR5RI8FMR0FLR2
RMVkOF0HMsR"CRl"5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GCRR5O8MFI08FR2CRslVRkH8GCRR5O8MFI08FR2RR=kGVHC58ROFR8IFM0R
82RkRVMHO0F"MRs"ClRR5D: R)qRp;sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-k-RVCHG8NR5RI8FMR0FLs2RCklRVCHG8NR5RI8FMR0Fj=2RRHkVGRC858NRF0IMFHRlMkHll,5Lj
22RkRVMHO0F"MRs"ClRR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GCRR5O8MFI0jFR2CRslVRkH8GCRR5O8MFI08FR2RR=kGVHC58ROFR8IFM0RMlHHllk5j8,2R2
RMVkOF0HMsR"CRl"5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8
;
R-R-RHkVGRC858NRF0IMF2RLR8lFRHkVGRC858NRF0IMF2RLRk=RVCHG8NR5RI8FMR0FLR2
RMVkOF0HMlR"FR8"5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GCRR5O8MFI08FR2FRl8VRkH8GCRR5O8MFI08FR2RR=kGVHC58ROFR8IFM0R
82RkRVMHO0F"MRl"F8RR5D: R)qRp;sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
R
R-k-RVCHG8NR5RI8FMR0FLl2RFk8RVCHG8NR5RI8FMR0Fj=2RRHkVGRC858NRF0IMFHRlMkHll,5Lj
22RkRVMHO0F"MRl"F8RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VRkH8GCRR5O8MFI0jFR2FRl8VRkH8GCRR5O8MFI08FR2RR=kGVHC58ROFR8IFM0RMlHHllk5j8,2R2
RMVkOF0HMlR"FR8"5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2+VR#H8GC58NRF0IMF2RLR#=RVCHG8+5N4FR8IFM0R
L2RkRVMHO0F"MR+5"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8OFR8IFM0RR82+VR#H8GC58ORF0IMF2R8R#=RVCHG8+5O4FR8IFM0R
82RkRVMHO0F"MR+5"RDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2+VR#H8GC58NRF0IMF2RjR#=RVCHG8+5N4FR8IFM0RMlHHllk5Lj,2R2
RMVkOF0HM+R""DR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RVCHG8R5O8MFI0jFR2RR+#GVHCO85RI8FMR0F8=2RRH#VG5C8OR+48MFI0lFRHlMHkjl5,282
VRRk0MOHRFM"R+"5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2-VR#H8GC58NRF0IMF2RLR#=RVCHG8+5N4FR8IFM0R
L2RkRVMHO0F"MR-5"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8OFR8IFM0RR82-VR#H8GC58ORF0IMF2R8R#=RVCHG8+5O4FR8IFM0R
82RkRVMHO0F"MR-5"RDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2-VR#H8GC58NRF0IMF2RjR#=RVCHG8+5N4FR8IFM0RMlHHllk5Lj,2R2
RMVkOF0HM-R""DR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RVCHG8R5O8MFI0jFR2RR-#GVHCO85RI8FMR0F8=2RRH#VG5C8OR+48MFI0lFRHlMHkjl5,282
VRRk0MOHRFM"R-"5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2*VR#H8GC58NRF0IMF2RLR#=RVCHG8N5.+84RF0IMFLR.2R
RVOkM0MHFR""*RR5D:hRz)m 1p7e _H#VG;C8R:sRRq) ps2RCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RVCHG8R5O8MFI08FR2RR*#GVHCO85RI8FMR0F8=2RRH#VG5C8.4O+RI8FMR0F.
82RkRVMHO0F"MR*5"RDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2*VR#H8GC58NRF0IMF2RjR#=RVCHG8N5.+84RF0IMF2RL
VRRk0MOHRFM"R*"5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8OFR8IFM0RRj2*VR#H8GC58ORF0IMF2R8R#=RVCHG8O5.+84RF0IMF2R8
VRRk0MOHRFM"R*"5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2/VR#H8GC58NRF0IMF2RLR#=RVCHG8-5NLR+48MFI0LFR-
N2RkRVMHO0F"MR/5"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8OFR8IFM0RR82/VR#H8GC58ORF0IMF2R8R#=RVCHG8-5O8R+48MFI08FR-
O2RkRVMHO0F"MR/5"RDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VG5C8NFR8IFM0RRL2/VR#H8GC58NRF0IMF2RjR#=RVCHG8+5N4FR8IFM0RNL-2R
RVOkM0MHFR""/RR5D:hRz)m 1p7e _H#VG;C8R:sRRaQh )t 2CRs0MksR)zh p1me_ 7#GVHC
8;
-RR-VR#H8GC58ORF0IMF2RjR#/RVCHG8R5O8MFI08FR2RR=#GVHCO85-48+RI8FMR0F-
O2RkRVMHO0F"MR/5"RDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

RR--#GVHC58RNFR8IFM0RRL2sRCl#GVHC58RNFR8IFM0RRL2=VR#H8GCRR5N8MFI0LFR2R
RVOkM0MHFRC"sl5"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VGRC858ORF0IMF2R8RlsCRH#VGRC858ORF0IMF2R8R#=RVCHG8OR5RI8FMR0F8R2
RMVkOF0HMsR"CRl"5:DRRq) ps;RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHC
8;
-RR-VR#H8GCRR5N8MFI0LFR2CRslVR#H8GCRR5N8MFI0jFR2RR=#GVHC58RNFR8IFM0RMlHHllk5jL,2R2
RMVkOF0HMsR"CRl"5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VGRC858ORF0IMF2RjRlsCRH#VGRC858ORF0IMF2R8R#=RVCHG8OR5RI8FMR0FlHHMl5kl82,j2R
RVOkM0MHFRC"sl5"RDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

RR--#GVHC58RNFR8IFM0RRL2lRF8#GVHC58RNFR8IFM0RRL2=VR#H8GCRR5N8MFI0LFR2R
RVOkM0MHFRF"l85"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VGRC858ORF0IMF2R8R8lFRH#VGRC858ORF0IMF2R8R#=RVCHG8OR5RI8FMR0F8R2
RMVkOF0HMlR"FR8"5:DRRq) ps;RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHC
8;
-RR-VR#H8GCRR5N8MFI0LFR2FRl8VR#H8GCRR5N8MFI0jFR2RR=#GVHC58RNFR8IFM0RMlHHllk5jL,2R2
RMVkOF0HMlR"FR8"5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsMz h)1emp #7_VCHG8
;
R-R-RH#VGRC858ORF0IMF2RjR8lFRH#VGRC858ORF0IMF2R8R#=RVCHG8OR5RI8FMR0FlHHMl5kl82,j2R
RVOkM0MHFRF"l85"RDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R

RR--a#EHRsPC#MHFRRFV8HHP8oCRH#PCRC0ERCk#sFRlsOCRFsM0FRD
RR--kGVHCN85RI8FMR0FL/2RRHkVG5C8OFR8IFM0RR82=VRkH8GC58N-RI8FMR0FL--O4R2
RMVkOF0HMHR8PCH8RR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8
RRRRMOF#M0N0FRsk_M8#D0$CRR:VCHG8F_sk_M8#D0$C$_0b:CR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRR:hzqa)RqpRRRRRRRRRRRRR:RR=HRVG_C8oskN8H_L0
#2RRRRskC0szMRh1) m pe7V_kH8GC;R

RR--a#EHRsPC#MHFRRFV8HHP8oCRH#PCRC0ERCk#sFRlsOCRFsM0FRD
RR--#GVHCN85RI8FMR0FL/2RRH#VG5C8OFR8IFM0RR82=VR#H8GC58N-+84RF0IMF-RLOR2
RMVkOF0HMHR8PCH8RR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8
RRRRMOF#M0N0FRsk_M8#D0$CRR:VCHG8F_sk_M8#D0$C$_0b:CR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRR:hzqa)RqpRRRRRRRRRRRRR:RR=HRVG_C8oskN8H_L0
#2RRRRskC0szMRh1) m pe7V_#H8GC;R

RR--a#ECCkRVMHO0FRM#skC0s4MR/RX
RR--4RR/kGVHCN85RI8FMR0FL=2RRHkVG5C8-8LRF0IMFNR--
42RkRVMHO0FsMRCbOHsNFOD
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRV:RH8GC_ksFM#8_0C$D_b0$C=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#Rh:Rq)azqRpRRRRRRRRRRRRRR=R:RGVHCo8_k8Ns_0LH#R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-4-RR#/RVCHG8R5N8MFI0LFR2RR=#GVHC-85LR+48MFI0-FRNR2
RMVkOF0HMCRsOsHbFDONRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR- R)vkRVMHO0FRM
RR--kGVHC58RNFR8IFM0RRL2sRClkGVHC58ROFR8IFM0R
82R-R-R=RRRHkVGRC85MlHHllk5ON,2FR8IFM0RMlHHllk58L,2R2
RMVkOF0HMCRslMNH8RCs5R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHC
8;RRRRO#FM00NMRksFM#8_0C$DRV:RH8GC_ksFM#8_0C$D_b0$C=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#Rh:Rq)azqRpRRRRRRRRRRRRRR=R:RGVHCo8_k8Ns_0LH#R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-#-RVCHG8NR5RI8FMR0FLs2RC#lRVCHG8OR5RI8FMR0F8R2
RR--RRR=#GVHC58RlHHMl5klN2,ORI8FMR0FlHHMl5klL2,82R
RVOkM0MHFRlsCN8HMC5sR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-FRl8kRVMHO0FRM
RR--kGVHC58RNFR8IFM0RRL2lRF8kGVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VRkH8GCRH5lMkHll,5NO82RF0IMFHRlMkHll,5LR282
VRRk0MOHRFMlkF8D5FR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7kGVHC
8;
-RR-VR#H8GCRR5N8MFI0LFR2FRl8VR#H8GCRR5O8MFI08FR2R
R-R-RRRRRRRR=#GVHC58ROFR8IFM0RMlHHllk5RL,8
22RkRVMHO0FlMRFD8kF
R5RRRRDs,RRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#RRRR:qRhaqz)pRRRRRRRRRRRRRRRRRRR:V=RH8GC_NoksL8_H20#
RRRR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RFusOkC8sVCRF0sRECF#RFIERCMC8MRNRO"NOkklDFN0sV"Rk0MOH3FM
-RR-8RN8N_OsRs$5HkVG5C8NFR8IFM0R,L2RHkVGRC858ORF0IMF2R82R
R-R-RRRRRR=RRRHkVGRC85GlNHllk5ON,2FR8IFM0RMlHHllk58L,2R2
RFbsOkC8sNCR8O8_N$ssRR5
RpRR,RR)RRR:HRMRz h)1emp k7_VCHG8R;
RORR_RHMRRR:HRMR1_a7ztpmQ
B;RRRRskC#D:0RR0FkR)zh p1me_ 7kGVHC
8;RRRROk_F0:RRR0FkR71a_mzpt2QB;R

RR--N_88OsNs$#R5VCHG8R5N8MFI0LFR2#,RVCHG8OR5RI8FMR0F8
22R-R-RRRRRRRRR#=RVCHG8lR5NlGHkNl5,RO28MFI0lFRHlMHkLl5,282
bRRsCFO8CksR8N8_sONs5$R
RRRRRp,)RRR:MRHRhRz)m 1p7e _H#VG;C8
RRRRHO_MRRR:MRHRaR17p_zmBtQ;R
RRCRs#0kDRF:Rkz0Rh1) m pe7V_#H8GC;R
RR_ROFRk0RF:Rk10Raz7_pQmtB
2;
-RR-OR1N#DCRC0ER#sCkRD0LN$RRIbFCFsRV3R.RHRW8R0EFHVRM0bkRI=RHE80RRFVFbk0kI0RH
0ER-R-RC0ERMLHNRs$bMFH0FRlP3C8
VRRk0MOHRFM#DONL$R5Rz:Rh1) m pe7V_kH8GC;RRh:hRQa  t)s2RCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM#DONL$R5Rz:Rh1) m pe7V_kH8GC;RRh:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMOR#NRDL5:$RR)zh p1me_ 7#GVHCR8;hRR:Q hat2 )R0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMOR#NRDL5:$RR)zh p1me_ 7#GVHCR8;hRR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _H#VG;C8
R
RVOkM0MHFR_Q#hNCo0CHPRs5NoRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp h
;
R-R-=========================================================================
==R-R-RlBFbHNs#RFMmsbCNs0F#R
R-=-==========================================================================R

RMVkOF0HM>R""5RRDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksRmAmph q;R
RVOkM0MHFR"">RDR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM"R<"R,5DR:sRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR<R"R5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM<R"=5"RDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksRmAmph q;R
RVOkM0MHFR="<"DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM"">=R,5DR:sRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR>R="5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM=R""5RRDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksRmAmph q;R
RVOkM0MHFR""=RDR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM""/=R,5DR:sRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR/R="5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp h
;
RkRVMHO0F"MR?R="R,5DR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"/R="5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR>"?"5RRDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R<"R,5DR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R="5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR="?"5RRDs,RRz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R>"R,5DR:sRR)zh p1me_ 7#GVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R">R="5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR<"?"5RRDs,RRz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;
VRRk0MOHRFM#_08lON0EDR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM#_08lON0EDR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
R
R-m-RPDCsF#N8RC0ERV8CN0kDRN"lGkHllN"RM"8RlHHMl"klRMVkOF0HMR

RMVkOF0HMNRlGkHllDR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMHRlMkHllDR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMNRlGkHllDR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMHRlMkHllDR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R--------------------------------------------------------------------------R-
RR--Q0MRECC#RlOFbCNsRMVkOF0HMN#RR0MNkDsNRRH#OPFMCCs08MRH0NFR
-RR-HRVGRC8bMFH0kRMlsLCRRFV0RECLMFk8"#RlHNGl5klDH'EojE,2FR8IFM0R
j"R-R--------------------------------------------------------------------------
-
RkRVMHO0F"MR=R"R5:DRR)zh p1me_ 7kGVHCR8;sRR:hzqa)2qpR0sCkRsMApmm ;qh
VRRk0MOHRFM""/=RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksRmAmph q;R
RVOkM0MHFR=">"DR5Rz:Rh1) m pe7V_kH8GC;RRs:qRhaqz)ps2RCs0kMmRAmqp hR;
RMVkOF0HM<R"=5"RDRR:z h)1emp k7_VCHG8s;RRh:Rq)azqRp2skC0sAMRm mpq
h;RkRVMHO0F"MR>R"R5:DRR)zh p1me_ 7kGVHCR8;sRR:hzqa)2qpR0sCkRsMApmm ;qh
VRRk0MOHRFM"R<"RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksRmAmph q;R

RMVkOF0HM=R""5RRDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR/R="5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM"">=RR5D:qRhaqz)ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksRmAmph q;R
RVOkM0MHFR="<"DR5Rh:Rq)azqRp;sRR:z h)1emp k7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM>R""5RRDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR<R"R5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh

RRRkRVMHO0F"MR?R="RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5Rz:Rh1) m pe7V_kH8GC;RRs:qRhaqz)ps2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR>"?=5"RDRR:z h)1emp k7_VCHG8s;RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R="5:DRR)zh p1me_ 7kGVHCR8;sRR:hzqa)2qpR0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R>"RR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5Rz:Rh1) m pe7V_kH8GC;RRs:qRhaqz)ps2RCs0kMaR17p_zmBtQ;R

RMVkOF0HM?R"=R"R5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?"/=RR5D:qRhaqz)ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5Rh:Rq)azqRp;sRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR<"?=5"RDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R">R"R5:DRRahqzp)q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R<"RR5D:qRhaqz)ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
R
RVOkM0MHFRGlNHllkRR5D:hRz)m 1p7e _HkVG;C8R:sRRahqzp)q2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0FlMRHlMHk5lRDRR:z h)1emp k7_VCHG8s;RRh:Rq)azq
p2RRRRskC0szMRh1) m pe7V_kH8GC;R
RVOkM0MHFRGlNHllkRR5D:qRhaqz)ps;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0FlMRHlMHk5lRDRR:hzqa);qpR:sRR)zh p1me_ 7kGVHC
82RRRRskC0szMRh1) m pe7V_kH8GC;R
R----------------------------------------------------------------------------
-RR-MRQRC0E#OCRFNlbsVCRk0MOH#FMRsNRCRNDHO#RFCMPs80CR0HMF
RNR-R-RGVHCb8RF0HMRlMkLRCsF0VRELCRF8kM#DR"'oEHER+48MFI0DFR'IDF"R
R----------------------------------------------------------------------------
R
RVOkM0MHFR""=RDR5Rz:Rh1) m pe7V_kH8GC;RRs: R)qRp2skC0sAMRm mpq
h;RkRVMHO0F"MR/R="5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksRmAmph q;R
RVOkM0MHFR=">"DR5Rz:Rh1) m pe7V_kH8GC;RRs: R)qRp2skC0sAMRm mpq
h;RkRVMHO0F"MR<R="5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksRmAmph q;R
RVOkM0MHFR"">RDR5Rz:Rh1) m pe7V_kH8GC;RRs: R)qRp2skC0sAMRm mpq
h;RkRVMHO0F"MR<R"R5:DRR)zh p1me_ 7kGVHCR8;sRR:)p q2CRs0MksRmAmph q;R

RMVkOF0HM=R""5RRDRR:)p q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM""/=RR5D: R)qRp;sRR:z h)1emp k7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM>R"=5"RDRR:)p q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM""<=RR5D: R)qRp;sRR:z h)1emp k7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM>R""5RRDRR:)p q;RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM"R<"RR5D: R)qRp;sRR:z h)1emp k7_VCHG8s2RCs0kMmRAmqp h
;
RkRVMHO0F"MR?R="RR5D:hRz)m 1p7e _HkVG;C8R:sRRq) ps2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR/"?=5"RDRR:z h)1emp k7_VCHG8s;RR):R 2qpR0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?">=RR5D:hRz)m 1p7e _HkVG;C8R:sRRq) ps2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR<"?=5"RDRR:z h)1emp k7_VCHG8s;RR):R 2qpR0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R>"RR5D:hRz)m 1p7e _HkVG;C8R:sRRq) ps2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR<"?"5RRDRR:z h)1emp k7_VCHG8s;RR):R 2qpR0sCkRsM1_a7ztpmQ
B;
VRRk0MOHRFM""?=RDR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"/R="5:DRRq) ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R="5:DRRq) ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R"R5:DRRq) ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
R
RVOkM0MHFRGlNHllkRR5D:hRz)m 1p7e _HkVG;C8R:sRRq) ps2RCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFMlHNGlRkl5:DRRq) ps;RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0FlMRHlMHk5lRDRR:z h)1emp k7_VCHG8s;RR):R 2qpR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMHRlMkHllDR5R):R ;qpR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R
R----------------------------------------------------------------------------
-RR-MRQRC0E#OCRFNlbsVCRk0MOH#FMRRNMHCM0oRCsHO#RFCMPs80CR0HMF
RNR-R-RGVHCb8RF0HMRlMkLRCsF0VRELCRF8kM#lR"NlGHkDl5'oEHE2,4RI8FMR0FjR"
R----------------------------------------------------------------------------R

RMVkOF0HM=R""5RRDRR:z h)1emp #7_VCHG8s;RRQ:Rhta  R)2skC0sAMRm mpq
h;RkRVMHO0F"MR/R="5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsMApmm ;qh
VRRk0MOHRFM"">=RR5D:hRz)m 1p7e _H#VG;C8R:sRRaQh )t 2CRs0MksRmAmph q;R
RVOkM0MHFR="<"DR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)s2RCs0kMmRAmqp hR;
RMVkOF0HM>R""5RRDRR:z h)1emp #7_VCHG8s;RRQ:Rhta  R)2skC0sAMRm mpq
h;RkRVMHO0F"MR<R"R5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsMApmm ;qh
R
RVOkM0MHFR""=RDR5RQ:Rhta  R);sRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM/R"=5"RDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR>R="5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM""<=RR5D:hRQa  t)s;RRz:Rh1) m pe7V_#H8GC2CRs0MksRmAmph q;R
RVOkM0MHFR"">RDR5RQ:Rhta  R);sRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp hR;
RMVkOF0HM<R""5RRDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0sAMRm mpq
h;
VRRk0MOHRFM""?=RDR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR/"?=5"RDRR:z h)1emp #7_VCHG8s;RRQ:Rhta  R)2skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R">R="5:DRR)zh p1me_ 7#GVHCR8;sRR:Q hat2 )R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?"<=RR5D:hRz)m 1p7e _H#VG;C8R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR<"?"5RRDRR:z h)1emp #7_VCHG8s;RRQ:Rhta  R)2skC0s1MRaz7_pQmtB
;
RkRVMHO0F"MR?R="RR5D:hRQa  t)s;RRz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5RQ:Rhta  R);sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR>"?=5"RDRR:Q hat; )R:sRR)zh p1me_ 7#GVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R="5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R>"RR5D:hRQa  t)s;RRz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5RQ:Rhta  R);sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R

RMVkOF0HMNRlGkHllDR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFMlHNGlRkl5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMHRlMkHllDR5Rz:Rh1) m pe7V_#H8GC;RRs:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFMlHHMlRkl5:DRRaQh )t ;RRs:hRz)m 1p7e _H#VG2C8
RRRR0sCkRsMz h)1emp #7_VCHG8R;
R----------------------------------------------------------------------------R
R-Q-RMER0CR#CObFlNRsCVOkM0MHF#RRNsDCNRRH#OPFMCCs08MRH0NFR
-RR-HRVGRC8bMFH0kRMlsLCRRFV0RECLMFk8"#RDH'Eo4E+RI8FMR0FDF'DIR"
R----------------------------------------------------------------------------R

RMVkOF0HM=R""5RRDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMApmm ;qh
VRRk0MOHRFM""/=RR5D:hRz)m 1p7e _H#VG;C8R:sRRq) ps2RCs0kMmRAmqp hR;
RMVkOF0HM>R"=5"RDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMApmm ;qh
VRRk0MOHRFM""<=RR5D:hRz)m 1p7e _H#VG;C8R:sRRq) ps2RCs0kMmRAmqp hR;
RMVkOF0HM>R""5RRDRR:z h)1emp #7_VCHG8s;RR):R 2qpR0sCkRsMApmm ;qh
VRRk0MOHRFM"R<"RR5D:hRz)m 1p7e _H#VG;C8R:sRRq) ps2RCs0kMmRAmqp h
;
RkRVMHO0F"MR=R"R5:DRRq) ps;RRz:Rh1) m pe7V_#H8GC2CRs0MksRmAmph q;R
RVOkM0MHFR="/"DR5R):R ;qpR:sRR)zh p1me_ 7#GVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR>R="5:DRRq) ps;RRz:Rh1) m pe7V_#H8GC2CRs0MksRmAmph q;R
RVOkM0MHFR="<"DR5R):R ;qpR:sRR)zh p1me_ 7#GVHCR82skC0sAMRm mpq
h;RkRVMHO0F"MR>R"R5:DRRq) ps;RRz:Rh1) m pe7V_#H8GC2CRs0MksRmAmph q;R
RVOkM0MHFR""<RDR5R):R ;qpR:sRR)zh p1me_ 7#GVHCR82skC0sAMRm mpq
h;
VRRk0MOHRFM""?=RDR5Rz:Rh1) m pe7V_#H8GC;RRs: R)qRp2skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"/R="5:DRR)zh p1me_ 7#GVHCR8;sRR:)p q2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5Rz:Rh1) m pe7V_#H8GC;RRs: R)qRp2skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R="5:DRR)zh p1me_ 7#GVHCR8;sRR:)p q2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5Rz:Rh1) m pe7V_#H8GC;RRs: R)qRp2skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R"R5:DRR)zh p1me_ 7#GVHCR8;sRR:)p q2CRs0MksR71a_mzpt;QB
R
RVOkM0MHFR="?"5RRDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?"/=RR5D: R)qRp;sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR>"?=5"RDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?"<=RR5D: R)qRp;sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFR>"?"5RRDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MR?R<"RR5D: R)qRp;sRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R

RMVkOF0HMNRlGkHllDR5Rz:Rh1) m pe7V_#H8GC;RRs: R)qRp2skC0szMRh1) m pe7V_#H8GC;R
RVOkM0MHFRGlNHllkRR5D: R)qRp;sRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFMlHHMlRkl5:DRR)zh p1me_ 7#GVHCR8;sRR:)p q2CRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0FlMRHlMHk5lRDRR:)p q;RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8R;
R=--=========================================================================R=
RR--1VEH0MRN8FR)0CN0RMwkOF0HM
#3R-R-R0hFCER0N#0RsNNRM#8RDNNRsMCRF00RE#CRNRlCN0#REACRQea_ mBa)CRPsF#HMR
R-=-==========================================================================R

RMVkOF0HM#R"DRD"5tq)Rz:Rh1) m pe7V_kH8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM"D#s"qR5):tRR)zh p1me_ 7kGVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMsR"FRD"5tq)Rz:Rh1) m pe7V_kH8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM"ssF"qR5):tRR)zh p1me_ 7kGVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HM#R"DRN"5tq)Rz:Rh1) m pe7V_kH8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM"N#s"qR5):tRR)zh p1me_ 7kGVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HM#R"DRD"5tq)Rz:Rh1) m pe7V_#H8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM"D#s"qR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMsR"FRD"5tq)Rz:Rh1) m pe7V_#H8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM"ssF"qR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HM#R"DRN"5tq)Rz:Rh1) m pe7V_#H8GC;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM"N#s"qR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HM]R1Q_wapa wRqR5):tRR)zh p1me_ 7kGVHCR8;BhmzaRR:hzqa)2qp
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HM]R1Q_wa)]QtaqR5):tRR)zh p1me_ 7kGVHCR8;BhmzaRR:hzqa)2qp
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HM]R1Q_wapa wRqR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:hzqa)2qp
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HM]R1Q_wa)]QtaqR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:hzqa)2qp
RRRR0sCkRsMz h)1emp #7_VCHG8
;
R-R--------------------------------------------------------------------------R-
RR--DHFoORNDVOkM0MHF#R
R----------------------------------------------------------------------------
R
RVOkM0MHFRF"M0R"R5RDRRRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM"8NM"5RRDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRFRs"RDR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMMR"N"M8R,5DR:sRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R
RVOkM0MHFRF"MsR"R5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVG;C8
VRRk0MOHRFM"sGF"5RRDs,RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRGsMF"DR5,RRs:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp k7_VCHG8R;
RMVkOF0HMMR"FR0"RR5DR:RRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R
RVOkM0MHFRM"N8R"R5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM""FsR5RRDs,RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRM8NM"DR5,RRs:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMMR"FRs"R,5DR:sRR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GC;R
RVOkM0MHFRF"GsR"R5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM"FGMs5"RDs,RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHC
8;
-RR-CReOs0FR8NMR8#0_FkDoRHOVOkM0MHF##,RNRlCNV#Rk0MOH#FMRRHMMCkls_HO#
08RkRVMHO0F"MRN"M8RDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRN"M8RDR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRFRs"RDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRFRs"RDR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRM8NM"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRM8NM"DR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRM"FsRDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRM"FsRDR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRG"FsRDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRG"FsRDR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRGsMF"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRGsMF"DR5Rz:Rh1) m pe7V_kH8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F"MRN"M8RDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRN"M8RDR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRFRs"RDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRFRs"RDR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRM8NM"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRM8NM"DR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRM"FsRDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRM"FsRDR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRG"FsRDR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRG"FsRDR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRGsMF"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RkRVMHO0F"MRGsMF"DR5Rz:Rh1) m pe7V_#H8GC;RRs:aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-CR)80kOHRFMFsbCNs0F##,RNRlCNM#RkslCH#O_0V8Rk0MOH#FM
VRRk0MOHRFM"8NM"5RRDRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFRN"MMR8"5:DRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HMFR"sR"RRR5D:hRz)m 1p7e _HkVG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRM"FsRDR5Rz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"sGF"5RRDRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFRM"GFRs"5:DRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HMNR"MR8"RR5D:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRM8NM"DR5Rz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""FsR5RRDRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQ;R
RVOkM0MHFRF"MsR"R5:DRR)zh p1me_ 7#GVHCR82skC0s1MRaz7_pQmtBR;
RMVkOF0HMGR"FRs"RR5D:hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRGsMF"DR5Rz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzpt;QB
R
R-s-RCs0kMN#RsDo'F4I-RRHVMRF0VMFk8R
RVOkM0MHFRMVH8C_DVF0l#50RNRso:hRz)m 1p7e _HkVG;C8R:$RR71a_mzpt2QB
RRRR0sCkRsMQ hat; )
VRRk0MOHRFMV8HM_VDC0#lF0NR5s:oRR)zh p1me_ 7#GVHCR8;$RR:1_a7ztpmQ
B2RRRRskC0sQMRhta  
);
-RR-CRs0Mks#sRNoH'Eo4E+RRHVMRF0VMFk8R
RVOkM0MHFRMVH8H_solE0FR#05oNsRz:Rh1) m pe7V_kH8GC;RR$:aR17p_zmBtQ2R
RRCRs0MksRaQh )t ;R
RVOkM0MHFRMVH8H_solE0FR#05oNsRz:Rh1) m pe7V_#H8GC;RR$:aR17p_zmBtQ2R
RRCRs0MksRaQh )t ;R

R=--=========================================================================R=
RR--R R)1 QZRMwkOF0HMR#
R=--=========================================================================R=
RR--sHC#xRC#0RECMLklC5sRDoNsCFsRslR#NCDDsR2
RR--aRECskC0s8MCR#sCkRD0IDHDRRLCkGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8GR2
RR--Q"VRsMFk80_#$"DCRRH#VCHG8F_sk,M8RC0EMER0CCRs#0kDRDIHDCRLRksFM88C3R
R-Q-RVER0C1RvAVRFRC0ERlsCN8HMCHsR#RRN"R4"qRh70RECpR1AF0VREkCRMksFM88CR#sCk
D0R-R-RRH#N4R''sRFRC0ERIDFCLsRHR0#F0VREsCRCHlNMs8CROHMDCk8R'NR40'RERCM0RECskC#DR0
RR--IDHDRRLCHsMOCCN#8$RLRC0ERN#lD#DC0CRsb#sCCNM0LRDCMLklCVsRF0sRERN00C$b3R
R-"-RFsPCVIDF_$#0DRC"ORNMLVCRH8GC_0#Nk0sNCsRFRGVHCI8_s3Nb
-RR-MRQR0#Nk0sNCFRl8RC,H0VREMCRkClLsPRFCDsVFRI#0MECRC0ERsDNo0C#R#bF#DHLCR
R-s-RCCbs#0CMNCLDRlMkLRCsHs#RCs0kM3C8RVRQRNIsbFRl8RC,0MECRC0ERbkbCLsRH
0#R-R-RRFV0RECMLklCNsRs0CRsOkMN80C3R
R
VRRk0MOHRFMsHC#x5CR
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-MRHb
k0RRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-H-RMo0CCbsRFHs0FRM
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;-RR-HR#xFCRVsRVNHO0FRM
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;
-RR-#R"H_xCs"C#RMVkOF0HMO#Rs0CNCER0CHR#xFCRVER0CkRF00bkRFVslER0CMRH8CHO#R
R-F-RVER0C#R"H_xCs"C#RbHMkR03RCaER0NOkRNDPkNDCVRFRH"#xsC_CR#"HM#RFk0R#3C8
VRRk0MOHRFMsHC#x5CR
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RsVFRx#HCMRFDR$
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;
-RR-FRh00CRERN0H"MRIbsN"FRl80CRE#CRHRoMLRH0HM#RFs0RCHbDOCN08R3Ra#EkRC0E
-RR-CRs#CHxRRFVNCRMoHN0PMCRkClLsNROMNREPNCRR#bFHP0HCCRs#0kDRRHMIbsNR8lFCR3
RMVkOF0HMCRs#CHxRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--HkMb0R
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )RRRRRRRRRRRR-H-RMo0CCbsRFHs0FRM
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;RRRRRRRRRRRRR--#CHxRRFVVOsN0MHF
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_#H8GC;R

RMVkOF0HMCRs#CHxRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--HkMb0R
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-V-RF#sRHRxCF$MD
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_#H8GC;R

R=--=========================================================================R=
RR--BPFMCHs#FwMRk0MOH#FM
-RR-===========================================================================
R
R-H-RMo0CC5sRMkN0s2NDRR0FkHM#o8MCRGVHCb8RF0HM3R
R-N-RslokC#M0RCNsRC0ERbkbCNsRMD8RFsICRkLFMR8#F0VREMCRkClLs0,RE
k#R-R-RHkVGRC858(RF0IMFdR-2=R<R_0FkGVHC58RH,M0RR(,-;d2
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:qRhaqz)pR;R-H-RMo0CCRs
RORRF0M#NRM0D0CV_8HMCRGRR:RRRaQh )t ;-RR-CRDVH0RMG8CRH5EoHERMG8C2R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hatR )RRRRRRRRRRRRRRRRR=R:RRj;RR--sEHo0MRH8
CGRRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
RVOkM0MHFR_0FkGVHC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRh:Rq)azqRp;RRRRRRRRR-RR-MRH0CCosR
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-V-RF#sRHRxCF$MD
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_kH8GC;R

RR--sDCNRR0FkHM#o8MCRGVHCb8RF0HM
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)qRp;RRRR-s-RC
NDRRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-D-RCRV0HCM8GER5HRoEHCM8GR2
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;-RR-HRsoRE0HCM8GR
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7kGVHC
8;
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)qRp;RRRR-s-RC
NDRRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RsVFRx#HCMRFDR$
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D;R
RRFROMN#0Mo0Rk8Ns_0LH#RRRRRR:hzqa)RqpRRRRRRRRRRRRRRRRR=R:RGVHCo8_k8Ns_0LH#R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-k-RMo#HMRC80kFRMo#HMRC8VCHG8FRbH
M0RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;RRRRRRRRRRRR-R-R#kMHCoM8R
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )R-R-RVDC0MRH8RCG5oEHEMRH82CG
RRRRMOF#M0N0HRso_E0HCM8GRRRRQ:Rhta  R)RRRRRRRRRRRRRRRRRRR:=jR;R-s-RH0oER8HMCRG
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7kGVHC
8;
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7R;RRRRRRRRRRR--kHM#o8MC
RRRRx#HCC_s#RRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-FRVsHR#xFCRM
D$RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-u-RCFsVsRl#NFROMsPC#MHF3kRRVCHG8NR5sso'NCMo2#RHR0sCkCsM8R
RVOkM0MHFR_0FkGVHC58R
RRRRoNsRz:Rh1) m pe7h_z1hQt R72RRRRRRRRRR--kHM#o8MC
RRRR0sCkRsMz h)1emp k7_VCHG8
;
R-R-R#kMHCoM8HRVGRC8bMFH0FR0R#kMHCoM8R
RVOkM0MHFR_0FkHM#o8MCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRRRRRRRR:hzqa);qpRRRRRRRRRRRR-D-RC0MoEVRFR0Fkb
k0RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _1zhQ th7
;
R-R-R#kMHCoM8HRVGRC8bMFH0FR0R#kMHCoM8R
RVOkM0MHFR_0FkHM#o8MCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;R-RR-HRVGRC8bMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7R;R-k-R#RC8VRFsDoCM0FERVkRF00bk
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7h_z1hQt 
7;
-RR-MRk#MHoCV8RH8GCRHbFM00RFCRsNRD
RMVkOF0HMFR0_NsCD
R5RRRRNRso:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM)p q;R

RR--kHM#o8MCRGVHCb8RF0HMRR0FHCM0o
CsRkRVMHO0F0MRFM_H0CCos
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksRahqzp)q;R

RR--QCM0oRCs0zFRh1) m pe7V_#H8GC
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRQa  t)R;RRR--HCM0o
CsRRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;RRR--D0CVR8HMC5GREEHoR8HMC
G2RRRRO#FM00NMRosHEH0_MG8CRRRR:hRQa  t)RRRRRRRRRRRRRRRRRRR:j=R;-RR-HRsoRE0HCM8GR
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$2DC
RRRR0sCkRsMz h)1emp #7_VCHG8
;
RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRaQh )t ;RRRRRRRRRRRRR--HCM0o
CsRRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RsVFRx#HCMRFDR$
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-CR)N0DRFVR#H8GC
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)qRp;RRRR-s-RC
NDRRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-D-RCRV0HCM8GER5HRoEHCM8GR2
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;-RR-HRsoRE0HCM8GR
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)qRp;RRRR-s-RC
NDRRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RsVFRx#HCMRFDR$
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D;R
RRFROMN#0Mo0Rk8Ns_0LH#RRRRRR:hzqa)RqpRRRRRRRRRRRRRRRRR=R:RGVHCo8_k8Ns_0LH#R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RHCoM8FR0RH#VG
C8RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 71hQt R7;RRRRRRRRRRRRR-R-Ro#HM
C8RRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-D-RCRV0HCM8GER5HRoEHCM8GR2
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t RRRRRRRRRRRRRRRRR:RR=;RjR-R-RosHEH0RMG8C
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_#H8GC;R

RMVkOF0HMFR0_H#VGRC85R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;R-#-RHCoM8R
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-V-RF#sRHRxCF$MD
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_#H8GC;R

RR--#MHoC08RFVR#H8GCRk5F00bkR#N#k8lCRR0FL#CRHRxCF#VRHCoM8MRHb2k0
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRso:hRz)m 1p7e _t1Qh2 7RRRRRRRRRRRR-#-RHCoM8R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-FRBMsPC#MHFRFVslVRkH8GCRR0F#GVHCR8
RMVkOF0HMFR0_H#VGRC85R
RRsRNoRR:z h)1emp k7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RHCoM8HRVGRC8bMFH0FR0Ro#HM
C8RkRVMHO0F0MRFH_#o8MCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRRRRRRRR:hzqa);qpRRRRRRRRRRRR-D-RC0MoEVRFR0Fkb
k0RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _t1Qh; 7
R
R-#-RHCoM8HRVGRC8bMFH0FR0Ro#HM
C8RkRVMHO0F0MRFH_#o8MCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;R-k-R#RC8VRFsDoCM0FERVkRF00bk
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7Q_1t7h ;R

RR--#MHoCV8RH8GCRHbFM00RFCRsNRD
RMVkOF0HMFR0_NsCD
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM)p q;R

RR--#MHoCV8RH8GCRHbFM00RFMRH0CCosR
RVOkM0MHFR_0FHCM0oRCs5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-V-RH8GCRHbFMH0RM0bk
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0sQMRhta  
);
-RR-CRAO#NkCVRFRC0ERHVNsRD$ObFlDNHO0RC8#HHxMsoRk#DCRRHM0RECVCHG8FRbH
M0R-R-RObN	CNo#ER0CR#CVOkM0MHF#sRNCsRbF8PHC08RFFROl0bkCER0CCRs#0kDRMsNo
C#R-R-RN GlCbD:R
R-#-RHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-#-RHNoMDVRk.RR:kGVHC58RcFR8IFM0R2-.;R
R-#-RHNoMDVRk4Dlk0.kVRk:RVCHG8kR5VCHG8H_Eo5ERd-,Rd',R*R',c-,R.82RF0IMFR
R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRkRRVCHG8F_DIdR5,dR-,*R''c,R,.R-2
2;R-R-R4kVl0kDkRV.<k=RV*4RR.kV;R
R-e-RN8DHRNOEs0NOC:s#R''+,-R''',R*R',',/'R''sRRFs'R)'5lsC2',RlF'RsvR''lR5F,82
-RR-RRRRRRRRRRRRRRRRRRR'R4'5OsCHFbsO2ND,NR''sRFR''qRL5N#R2,'RM'F'sRh5'RksMN$2R-
VRRk0MOHRFMkGVHCE8_HRoE5VDC0M_H8,CGRosHEH0_MG8CR:RRRaQh )t ;R
RRRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMRRRRRRRRRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMC,G.RosHEH0_MG8C.RR:Q hatR )R=R:R
j2RRRRskC0sQMRhta  
);RRR
RMVkOF0HMVRkH8GC_IDFRC5DVH0_MG8C,HRso_E0HCM8GRRR:hRQa  t)R;
RRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMRRRRRRRRRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GR.,sEHo0M_H8.CGRQ:Rhta  R)RRR:=jR2
RsRRCs0kMhRQa  t)R;
RR
RVOkM0MHFRH#VG_C8EEHoRC5DVH0_MG8C,HRso_E0HCM8GRRR:hRQa  t)R;
RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRRRRRRRRRRRRRRRRRB:R]qq)B)a RR:=';X'
RRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8.CG,HRso_E0HCM8G:.RRaQh )t R:RR=2Rj
RRRR0sCkRsMQ hat; )

RRRkRVMHO0F#MRVCHG8F_DIDR5C_V0HCM8Gs,RH0oE_8HMCRGRRQ:Rhta  
);RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRRRRRRRRRRRRRRRRRB:R]qq)B)a RR:=';X'
RRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMC,G.RosHEH0_MG8C.RR:Q hatR )R=R:R
j2RRRRskC0sQMRhta  
);
-RR-NR1lNCR#LRNF,PCR0LkRHk#M0oRE"CR#CHx_#sC"MRHbRk0F$MDRsVFRC0EHssRNCMo#R:
RR--#MHoNkDRVk4lDV0k.RR:kGVHC58RkGVHCE8_HRoE54kV,*R''k,RVR.28MFI0RF
RR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRkGVHCD8_F5IRk,V4R''*,VRk.;22
-RR-VRk4Dlk0.kVRR<=kRV4*VRk.R;
RR--
VRRk0MOHRFMkGVHCE8_HRoE5x#HCC_s#:RRR)zh p1me_ 7kGVHC
8;RRRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRRRRRHR#xsC_CR#.:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMQ hat; )

RRRkRVMHO0FkMRVCHG8F_DI#R5H_xCsRC#Rz:Rh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRRRRRRCFbsHN0F:MRRqB])aqB :)R=XR''R;
RRRRRRRRRRRRRRRRRRRRRHR#xsC_CR#.:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMQ hat; )

RRRkRVMHO0F#MRVCHG8H_Eo5ER#CHx_#sCRRR:z h)1emp #7_VCHG8R;
RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRB:R]qq)B)a RR:=';X'
RRRRRRRRRRRRRRRRRRRRRRRRx#HCC_s#:.RR)zh p1me_ 7#GVHC
82RRRRskC0sQMRhta  
);RRR
RMVkOF0HMVR#H8GC_IDFRH5#xsC_CR#R:hRz)m 1p7e _H#VG;C8
RRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRRRRRx#HCC_s#:.RR)zh p1me_ 7#GVHC
82RRRRskC0sQMRhta  
);
-RR-kRbs#bFCs:RCs0kMN#RR0#Nk0sNCM8RkClLsR
RVOkM0MHFR0#Nk0sNC
R5RRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC;R

RR--bbksF:#CR0sCk#sMR#NRNs0kN80CRlMkL
CsRkRVMHO0F#MRNs0kNR0C5R
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t ;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
VRRk0MOHRFM#kN0sCN0RR5
R#RRH_xCsRC#:hRz)m 1p7e _HkVG2C8RRRRR-RR-MRFD0$RE#CRHRxCF0VRERH#Hk#R#
C8RRRRskC0szMRh1) m pe7V_kH8GC;R

RMVkOF0HMNR#0Nks05CR
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2RRRRRRR--F$MDRC0ERx#HCVRFRH0E##RHRCk#8R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-===========================================================================
-RR-sRaNDM#NF0HMkRwMHO0F
M#R-R-=========================================================================
==
-RR-NRlbl#RC-0NDHFoORNDPkNDCR#
RMVkOF0HMFR0_Rj45R
RRRR#RRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0XuvqR1:Raz7_pQmtB=R:R''j2-RR-NRvbRRG0RF
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-l-RNRb#lNC0-oDFHDONRDPNk
C#RkRVMHO0F0MRF4_jRR5
R#RRRRRRRRRRRRRRRz:Rh1) m pe7V_#H8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRO#FM00NMRqXvuRR:1_a7ztpmQ:BR=jR''R2R-v-RNGbRR
0FRRRRskC0szMRh1) m pe7V_#H8GC;R

RMVkOF0HM#RQ_RXRRNR5s:oRR)zh p1me_ 7kGVHCR82skC0sAMRm mpq
h;RkRVMHO0FQMR#R_XR5RRNRso:hRz)m 1p7e _H#VG2C8R0sCkRsMApmm ;qh
VRRk0MOHRFM0XF_jR4R5oNsRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F0MRFj_X45RRNRso:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8R;
RMVkOF0HMFR0_4XjZNR5s:oRR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GC;R
RVOkM0MHFR_0FXZj4Rs5NoRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VG;C8
VRRk0MOHRFM0zF_XRj45oNsRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHC
8;RkRVMHO0F0MRFX_zj54RNRso:hRz)m 1p7e _H#VG2C8R0sCkRsMz h)1emp #7_VCHG8
;
R-R-Rs#0NEHo0CRPOs0FRMOFP#CsHRFMs0FkH#MC,CRMC88CRsVFRM#$0#ECH
#3R-R-RCaE#VCRk0MOH#FMRCNsRsECCFR#RN0E0RRN#_08DHFoOC_POs0FRMONR
LCR-R-RMOFP0CsC08RFMRN8sRVF#lRVCHG8MRN8VRkH8GC3hRRFR0C00ENRk$FRMON
-RR-FRM0FROMsPC0ER0CR#CP0COFRs#LNCOkR#CF0VREsCHRoMCNP0HCMRH83CG

RRRkRVMHO0F0MRFD_#P
R5RRRRNRso:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRR-V-RH8GCRHbFMP0RCFO0sR
RRCRs0MksR71a_tpmQeB_ mBa)R;
RHNDN0#RF0_18opFHCOeOs0FRRH#0#F_DrPRz h)1emp k7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR17m_pt_QBea Bm;)9
NRRD#HNR_0F1_08pHFoOC_eOs0FRRH#0#F_DrPRz h)1emp k7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM1_a7pQmtB _eB)am9
;
RkRVMHO0F0MRFD_#P
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-V-RH8GCRHbFMP0RCFO0sR
RRCRs0MksR71a_tpmQeB_ mBa)R;
RHNDN0#RF0_18opFHCOeOs0FRRH#0#F_DrPRz h)1emp #7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMaR17m_pt_QBea Bm;)9
NRRD#HNR_0F1_08pHFoOC_eOs0FRRH#0#F_DrPRz h)1emp #7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsM1_a7pQmtB _eB)am9
;
RkRVMHO0F0MRFk_#D5PR
RRRRoNsRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRRR--VCHG8FRbHRM0P0COFRs
RsRRCs0kMaR17p_zmBtQ_Be a;m)
NRRD#HNR_0F1z08pHFoOOeC0RFsH0#RFk_#DrPRz h)1emp k7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0s1MRaz7_pQmtB _eB)am9R;
RHNDN0#RF0_18p_zFOoH_OeC0RFsH0#RFk_#DrPRz h)1emp k7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR71a_mzpt_QBea Bm;)9
R
RVOkM0MHFR_0F#PkDRR5
RNRRs:oRR)zh p1me_ 7#GVHCR82RRRRRRRRR-RR-HRVGRC8bMFH0CRPOs0F
RRRR0sCkRsM1_a7ztpmQeB_ mBa)R;
RHNDN0#RF0_18FzpoeHOCFO0s#RHR_0F#PkDRhrz)m 1p7e _H#VG
C8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR71a_mzpt_QBea Bm;)9
NRRD#HNR_0F1_08zopFHeO_CFO0s#RHR_0F#PkDRhrz)m 1p7e _H#VG
C8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0s1MRaz7_pQmtB _eB)am9
;
RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRR:aR17p_zmBtQ_Be a;m)R-R-RH#EV80CROPC0
FsRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC;R

RMVkOF0HMFR0_HkVGRC85R
RRsRNoRRRR:RRR71a_mzpt_QBea BmR);RRRRR-R-RH#EV80CROPC0
FsRRRR#CHx_#sCRz:Rh1) m pe7V_kH8GC2RRRRRRR-V-RF#sRHRxCF$MD
RRRR0sCkRsMz h)1emp k7_VCHG8
;
RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRR:aR17p_zmBtQ_Be a;m)R-R-RH#EV80CROPC0
FsRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC;R

RMVkOF0HMFR0_H#VGRC85R
RRsRNoRRRR:RRR71a_mzpt_QBea BmR);RRRRR-R-RH#EV80CROPC0
FsRRRR#CHx_#sCRz:Rh1) m pe7V_#H8GC2RRRRRRR-V-RF#sRHRxCF$MD
RRRR0sCkRsMz h)1emp #7_VCHG8
;
R-R-RRq#NFROM#OC#MHFRR0F0#EFCERIF#RkCRRNobsNENHOD1R7uMRCPFHsMMlC0R,
RR--0#ECCkRVMHO0FRM#0CN	RsbNN0lCCRs#H0MRECF#RF0FDV#RFNsl0MRN8sROCCN0
-RR-HRVGRC8bMFH0kRMlsLC#R3Ra#ECCkRVMHO0FRM#NRsC8HC#o8MCRR0FOPFMCRs0VlsF
-RR-RRN#_08DHFoOC_POs0FRR0F0RECep]7RGVHCb8RF0HMRsVFlRN0kM#HoER0CFROMMPC0MHF#R
R-F-RVER0CR#Cb	NON#oC3QRRMRRNbCksR7e]pMRCPFHsMMlC0FR$kER#F8kDRCk#RC0E
-RR-0R"FV_kH8GC"MRN80R"FV_#H8GC"FRskM0HC
#3
-RR-MRk#MHoCV8RH8GCRHbFMR0
RMVkOF0HMFR0_HzwG
R5RRRRNRsoRRRRR1:Raz7_pQmtB _eB)am;R
RRHRI8R0ER:RRRahqzp)q;RRRRRRRRRRRRRRRR-R-R8IH0FERVCRPOs0F
RRRRNVsOF0HMRR:hzqa)2qpRRRRRRRRRRRRRRRRRR--I0H8EVRFRNVsOF0HMR
RRCRs0MksR)zh p1me_ 7kGVHC
8;
-RR-HR#o8MCRGVHCb8RF0HM
VRRk0MOHRFM01F_wRHG5R
RRsRNoRRRR:RRR71a_mzpt_QBea Bm
);RRRRI0H8ERRRRh:Rq)azqRp;RRRRRRRRRRRRRRRR-I-RHE80RRFVP0COFRs
RVRRs0NOHRFM:qRhaqz)pR2RRRRRRRRRRRRRR-RR-HRI8R0EFVVRs0NOH
FMRRRRskC0szMRh1) m pe7V_#H8GC;R

RR--V8HMHRMo0RECLMFk8F#RVRRNMLklCRs3RCaE#VCRk0MOH#FMRMONRRLCk8#CR	DHCER0H
#:R-R-Ro#HMRNDGRGG:VRkH8GCRR5(8MFI0-FRd
2;R-R-RR--WOEHE#RHRC0ERl#NC#RNRV"kH8GCRw5zHEG_HRoE5,44d82RF0IMFwRzHDG_F4I542,d2R"
RR--#MHoN$DR$:$RRHkVGRC85HzwGH_Eo5ER4R4,d",R+R",4R4,dR2
RR--RRRRRRRRRRRRRFR8IFM0RHzwGF_DI454,,RdR""+,4R4,2Rd2R;
RR--WsECC4R"4H"R#ER0CHRI8R0EFGVRG5GRG'GGDoCM0,E2
-RR-MRN8RRdH0#REDCRFsICRkLFM58RNRL#5GGG'IDF2R2
RR--QNMRRsbkC]Re7CpRMsPHFCMlMk0R#"CRkGVHCE8_H"oER8NMRV"kH8GC_IDF"R
R
VRRk0MOHRFMzGwH_oEHEIR5HE80,sRVNHO0FRMRRh:Rq)azq
p;RRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRRHRI8.0E,sRVNHO0FRM.:qRhaqz)pRRR:j=R2R
RRCRs0MksRaQh )t ;R
R
VRRk0MOHRFMzGwH_IDFRH5I8,0ERNVsOF0HMRRR:qRhaqz)pR;
RRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRRRRRRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRIRRHE80.V,Rs0NOH.FMRh:Rq)azqRpRRR:=jR2
RsRRCs0kMhRQa  t)
;
R-R-Rl1NC#RNRFNLPLCRkV0RF#sRHCoM8HRVGRC8bMFH0R3RhCF0RN0E0ER0CHRI8
0ER-R-RRFVNHR#o8MCRGVHCb8RF0HMRlMkLRCsHFoMsRC#0REC#MHoR0LH,ER0kR#
RR--I0H8ERR=#GGG'MDCo-0E4R
R
VRRk0MOHRFM1GwH_oEHEIR5HE80,sRVNHO0FRMRRh:Rq)azq
p;RRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRRHRI8.0E,sRVNHO0FRM.:qRhaqz)pRRR:j=R2R
RRCRs0MksRaQh )t ;R
R
VRRk0MOHRFM1GwH_IDFRH5I8,0ERNVsOF0HMRRR:qRhaqz)pR;
RRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRRRRRRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRIRRHE80.V,Rs0NOH.FMRh:Rq)azqRpRRR:=jR2
RsRRCs0kMhRQa  t)
;
R-R-=========================================================================
==R-R-Rs#0HRMoNRM800CGHwFRk0MOH#FM
-RR-===========================================================================
-
-bosNl#NR$EM0C##H_VFV
R--s_0D#0$MEHC##VRFVR

RR--bbksF:#CRHIs0RC#VCHG8FRbHRM0HFM0RDNRH
MCRsRbF8OCkRsCWa)Q 
R5RRRRpRRRRRRRRRR:HkMF0QRphR ;RRRRRRRRRRRRR-R-RbHMkD0RH
MCRRRRezqp RRRRRR:HRMRRhRz)m 1p7e _HkVG;C8R-R-RGVHCb8RF0HMRbHMkR0
RKRRzQ1aw7Q RH:RMRRRR71Q :RR=HRso;E0
RRRR wQpR7RR:RRRRHMRWRRQ]7aRR:=j
2;
-RR-kRbs#bFCI:RsCH0#HRVGRC8bMFH0MRH0NFRRMDHCR
RbOsFCs8kC)RWQRa 5R
RRRRpRRRRRRRR:MRHFRk0p Qh;RRRRRRRRRRRRRRR-H-RM0bkRMDHCR
RRqRepRz RRRR:MRHRRRRz h)1emp #7_VCHG8R;R-V-RH8GCRHbFMH0RM0bk
RRRR1KzaQQw :7RRRHMR1RRQR7 RR:=sEHo0R;
RwRRQ7 pRRRRRH:RMRRRR7WQa:]R=2Rj;R

RFbsOkC8s)CR 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_kH8GC2
;
RsRbF8OCkRsC)7 q5RpRR:RRRFHMkp0RQ;h 
RRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp k7_VCHG8R;
RRRRRRRRRRRRRRRRt7mmRRR:FRk0RmRAmqp h
2;
bRRsCFO8CksRq) 7R5pRRRR:MRHFRk0p Qh;R
RRRRRRRRRRRRRReRRq pzRF:RkR0RR)zh p1me_ 7#GVHC;82
R
RbOsFCs8kC R)qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRezqp RR:FRk0RhRz)m 1p7e _H#VG;C8
RRRRRRRRRRRRRRRRmRtmR7R:kRF0RRRApmm 2qh;R

RHNDNL#RI0sHC#RHRQW)ar Rp Qh,hRz)m 1p7e _HkVG,C8R71Q I,RHE809R;
RHNDNL#RI0sHC#RHRQW)ar Rp Qh,hRz)m 1p7e _H#VG,C8R71Q I,RHE809R;
RHNDNL#Rs8CNRRH#)7 qRQrphR ,z h)1emp k7_VCHG8
9;RDRNHRN#LNsC8#RHRq) 7pRrQ,h R)zh p1me_ 7kGVHCR8,Apmm 9qh;R
RNNDH#sRLCRN8H)#R Rq7rhpQ z,Rh1) m pe7V_#H8GC9R;
RHNDNL#Rs8CNRRH#)7 qRQrphR ,z h)1emp #7_VCHG8A,Rm mpq;h9
NRRD#HNRhAQq_)YWa)Q #RHRQW)ar Rp Qh,hRz)m 1p7e _HkVG,C8R71Q I,RHE809R;
RHNDNA#RQ)hqY)_WQRa HW#R) QaRQrphR ,z h)1emp #7_VCHG81,RQ,7 R8IH0;E9
NRRD#HNRhAQq_)Y)7 qRRH#)7 qRQrphR ,z h)1emp k7_VCHG8A,Rm mpq;h9
NRRD#HNRhAQq_)Y)7 qRRH#)7 qRQrphR ,z h)1emp k7_VCHG8
9;RDRNHRN#AqQh))Y_ Rq7H)#R Rq7rhpQ z,Rh1) m pe7V_#H8GC,mRAmqp h
9;RDRNHRN#AqQh))Y_ Rq7H)#R Rq7rhpQ z,Rh1) m pe7V_#H8GC9
;
R-R-R0FONsDRCRN8NRM8I0sHCR
RbOsFCs8kCWRm) QaRR5
RpRRRRRRRRRRRH:RM0FkRhpQ R;RRRRRRRRRRRRRRR--HkMb0HRDMRC
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7kGVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2
;
RsRbF8OCkRsCmQW)a5 R
RRRRRpRRRRRR:RRRFHMkp0RQ;h RRRRRRRRRRRRR-RR-MRHbRk0DCHM
RRRRpeqzR RR:RRRRHMRzRRh1) m pe7V_#H8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRKaz1Q wQ7RR:HRMRRQR17R R:s=RH0oE;R
RRQRw Rp7RRRR:MRHRRRRWaQ7]=R:R;j2
R
RbOsFCs8kC)Rm 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp k7_VCHG8
2;
bRRsCFO8CksR m)qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRt7mmRRR:FRk0RmRAmqp h
2;
bRRsCFO8CksR m)qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_#H8GC2
;
RsRbF8OCkRsCmq) 7R5pRRRR:MRHFRk0p Qh;R
RRRRRRRRRRRRRRRRRezqp RR:FRk0RhRz)m 1p7e _H#VG;C8
RRRRRRRRRRRRRRRRtRRmRm7RF:RkR0RRmAmph q2R;
RHNDNm#RBpaq_q) 7#RHR m)qr7Rp Qh,hRz)m 1p7e _HkVG,C8RmAmph q9R;
RHNDNm#RBpaq_q) 7#RHR m)qr7Rp Qh,hRz)m 1p7e _HkVG9C8;R
RNNDH#BRma_qp)7 qRRH#mq) 7pRrQ,h R)zh p1me_ 7#GVHCR8,Apmm 9qh;R
RNNDH#BRma_qp)7 qRRH#mq) 7pRrQ,h R)zh p1me_ 7#GVHC;89
NRRD#HNRamBqWp_) QaRRH#mQW)ar Rp Qh,hRz)m 1p7e _HkVG,C8R71Q W,RQ]7a9R;
RHNDNm#RBpaq_QW)aH R#WRm) QaRQrphR ,z h)1emp #7_VCHG81,RQ,7 R7WQa;]9
R
R-E-RCsGRCRN8NRM8I0sHCR
RbOsFCs8kCWR]) QaRR5
RpRRRRRRRRRRRH:RM0FkRhpQ R;RRRRRRRRRRRRRRR--HkMb0HRDMRC
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7kGVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2
;
R-R-RsbkbCF#:sRIH#0CRGVHCb8RF0HMR0HMFRRNDCHM
bRRsCFO8CksR)]WQRa 5R
RRRRpRRRRRRRR:MRHFRk0p Qh;RRRRRRRRRRRRRRR-H-RM0bkRMDHCR
RRqRepRz RRRR:MRHRRRRz h)1emp #7_VCHG8R;R-V-RH8GCRHbFMH0RM0bk
RRRR1KzaQQw :7RRRHMR1RRQR7 RR:=sEHo0R;
RwRRQ7 pRRRRRH:RMRRRR7WQa:]R=2Rj;R

RFbsOkC8s]CR)7 q5RpRR:RRRFHMkp0RQ;h 
RRRRRRRRRRRRRRRReRRq pzRF:RkR0RR)zh p1me_ 7kGVHC;82
R
RbOsFCs8kC)R] 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp k7_VCHG8R;
RRRRRRRRRRRRRRRRRmtm7:RRR0FkRARRm mpq;h2
R
RbOsFCs8kC)R] 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp #7_VCHG8
2;
bRRsCFO8CksR ])qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_#H8GC;R
RRRRRRRRRRRRRRRRRt7mmRRR:FRk0RmRAmqp h
2;RDRNHRN#]_ X)7 qRRH#]q) 7pRrQ,h R)zh p1me_ 7kGVHCR8,Apmm 9qh;R
RNNDH# R]X _)qH7R#)R] Rq7rhpQ z,Rh1) m pe7V_#H8GC,mRAmqp h
9;RDRNHRN#]_ X)7 qRRH#]q) 7pRrQ,h R)zh p1me_ 7kGVHC;89
NRRD#HNRX] _q) 7#RHR ])qr7Rp Qh,hRz)m 1p7e _H#VG9C8;R
RNNDH# R]X)_WQRa H]#RWa)Q pRrQ,h R)zh p1me_ 7kGVHCR8,1 Q7,QRW79a];R
RNNDH# R]X)_WQRa H]#RWa)Q pRrQ,h R)zh p1me_ 7#GVHCR8,1 Q7,QRW79a];R

RR--skC0sRM#N0R#soHM,#RkCDVkRsVF:R
R-N-R#s#C0GR5R$=R2CRsb0FsRs"CsRFsVMFk8RR"&FR0_s#0H5MoG#2RCsPCHR0$CFsssR;
RMVkOF0HMFR0_s#0HRMo5DPNk:CRR)zh p1me_ 7kGVHCR82skC0s1MRah)Qt
;
RDRNHRN#0LF_#H0sMHoR#FR0_s#0HRMor)zh p1me_ 7kGVHCs8RCs0kMaR1)tQh9R;
RHNDNa#RmQ_AhYq)_)1aQRhtHa#Rma_1)tQhRhrz)m 1p7e _HkVGRC8skC0s1MRah)Qt
9;
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:z h)1emp k7_VCHG8s2RCs0kMaR1)tQh;R
RNNDH#mRa_amBq1p_ah)Qt#RHR_amm)1aQRhtr)zh p1me_ 7kGVHCs8RCs0kMaR1)tQh9
;
RkRVMHO0F0MRF#_E0MsHoPR5NCDkRz:Rh1) m pe7V_kH8GC2CRs0MksR)1aQ;ht
NRRD#HNR_am]_ X1Qa)hHtR#mRa_a]1)tQhRhrz)m 1p7e _HkVGRC8skC0s1MRah)Qt
9;
VRRk0MOHRFM0#F_0MsHoPR5NCDkRz:Rh1) m pe7V_#H8GC2CRs0MksR)1aQ;ht
NRRD#HNR_0FLs#0HRMoH0#RF0_#soHMRhrz)m 1p7e _H#VGRC8skC0s1MRah)Qt
9;RDRNHRN#aAm_Q)hqYa_1)tQhRRH#a1m_ah)QtzRrh1) m pe7V_#H8GCR0sCkRsM1Qa)h;t9
R
RVOkM0MHFR_0FFs#0HRMo5DPNk:CRR)zh p1me_ 7#GVHCR82skC0s1MRah)QtR;
RHNDNa#RmB_ma_qp1Qa)hHtR#mRa_am1)tQhRhrz)m 1p7e _H#VGRC8skC0s1MRah)Qt
9;
VRRk0MOHRFM0EF_#H0sM5oRPkNDCRR:z h)1emp #7_VCHG8s2RCs0kMaR1)tQh;R
RNNDH#mRa_X] _)1aQRhtHa#Rm1_]ah)QtzRrh1) m pe7V_#H8GCR0sCkRsM1Qa)h;t9
R
R-w-RsRFl#H0sMVoRk0MOH#FMRDNDF$IRF0kRFFROMsPC0RRN#H0sMHoRMR0FNHRVG
C8R-R-RHbFMM0RkClLsR3R lGNb:DC
-RR-#RRHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-R-RkRV4<V=Rs_Fl#H0sM5oR"4j4jj34jR",k'V4EEHo,VRk4F'DIR2;-n-R3R6
RR--aREC"R3"HF#RbF0HMRNDH0MRERH##0$MNRG,ECFIPRCsHC0RG0H#R8NMR
H#R-R-RRHM0RECIMsFoFRDOHN0FNMRMsRCsRFsHb#RskF8O3C8RPRmCDsVFIIRH
DDR-R-R#sCkRD0H#MRNs0kNF0HMR3
RR
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoRRRRRRRRRRRRR:aR1)tQh;RRRR-RR-HRLM$NsRs#0H
MoRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC;R
RNNDH#sRVFLl_#H0sMHoR#sRVF#l_0MsHo1Rrah)QtQ,Rhta  R),Q hat
 )RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp k7_VCHG8
9;RDRNHRN#VlsF_MLHN_s$#H0sMHoR#sRVF#l_0MsHo1Rrah)QtQ,Rhta  R),Q hat
 )RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _HkVG9C8;R

RR--mNO0DMRN8CREGFROMsPC#MHF#FRIsN	R#FRVDIDF#R:
RR--kRV4<V=Rs_FlEs#0HRMo53"nUR",d-,RdR2;-n-R356RL0F0FxlRC#sFRF8sb8bC2R
R-k-RV<4R=sRVFFl_#H0sM5oR"3jncR",d-,RdR2;-n-R356R0RFbxFCs#sR8FCbb8R2
RR
RVOkM0MHFRFVsl#_F0MsHo
R5RRRRFs#0HRMoRRRRRRRRRRRRR1:Rah)QtR;RRRRR-m-ROD0NRs#0H
MoRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC;R
RNNDH#sRVFFl_OD0N_s#0HRMoHV#Rs_FlFs#0HRMor)1aQ,htRaQh )t ,hRQa  t)R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp k7_VCHG8
9;
VRRk0MOHRFMVlsF_0E#soHMRR5
RERR#H0sMRoRRRRRRRRRRRRR:aR1)tQh;RRRR-RR-CREG0R#soHM
RRRRMOF#M0N0CRDVH0_MG8CRRR:Q hat; )
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hat2 )
RRRR0sCkRsMz h)1emp k7_VCHG8R;
RHNDNV#Rs_FlE_CG#H0sMHoR#sRVFEl_#H0sMroR1Qa)hRt,Q hat, )RaQh )t 
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7kGVHC;89
R
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoRRRRRRRRRRRRR:aR1)tQh;RRRR-RR-HRLM$NsRs#0H
MoRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC;R
RNNDH#sRVFLl_#H0sMHoR#sRVF#l_0MsHo1Rrah)QtQ,Rhta  R),Q hat
 )RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp #7_VCHG8
9;RDRNHRN#VlsF_MLHN_s$#H0sMHoR#sRVF#l_0MsHo1Rrah)QtQ,Rhta  R),Q hat
 )RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _H#VG9C8;R

RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRRRRRRRRRRRRRR:1Qa)hRt;RRRRRR--mNO0D0R#soHM
RRRRMOF#M0N0CRDVH0_MG8CRRR:Q hat; )
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R;
RHNDNV#Rs_FlFNO0D0_#soHMRRH#VlsF_0F#soHMRar1)tQh,hRQa  t)Q,Rhta  R)
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7#GVHC;89
R
RVOkM0MHFRFVsl#_E0MsHo
R5RRRREs#0HRMoRRRRRRRRRRRRR1:Rah)QtR;RRRRR-E-RC#GR0MsHoR
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t ;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RDRNHRN#VlsF_GEC_s#0HRMoHV#Rs_FlEs#0HRMor)1aQ,htRaQh )t ,hRQa  t)R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _H#VG9C8;R

RR--1CNlRRN#NPLFC",R#CHx_#sC"#RHRCk#8FRVs0RH's#RNCMoRDFM$R3
RMVkOF0HMsRVF#l_0MsHo
R5RRRRLs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-L-RHsMN$0R#soHM
RRRRx#HCC_s#RR:z h)1emp k7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
NRRD#HNRFVsl#_L0MsHo#RHRFVsl0_#soHMRar1)tQh,hRz)m 1p7e _HkVG
C8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp k7_VCHG8
9;RDRNHRN#VlsF_MLHN_s$#H0sMHoR#sRVF#l_0MsHo1Rrah)Qtz,Rh1) m pe7V_kH8GC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0szMRh1) m pe7V_kH8GC9
;
RkRVMHO0FVMRs_FlFs#0HRMo5R
RR#RF0MsHo:RRR)1aQ;htRRRRRRRRRRRRRRRRR-R-R0mON#DR0MsHoR
RRHR#xsC_C:#RR)zh p1me_ 7kGVHC
82RRRRskC0szMRh1) m pe7V_kH8GC;R
RNNDH#sRVFFl_OD0N_s#0HRMoHV#Rs_FlFs#0HRMor)1aQ,htR)zh p1me_ 7kGVHCR8
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7kGVHC;89
R
RVOkM0MHFRFVsl#_E0MsHo
R5RRRREs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-E-RC#GR0MsHoR
RRHR#xsC_C:#RR)zh p1me_ 7kGVHC
82RRRRskC0szMRh1) m pe7V_kH8GC;R
RNNDH#sRVFEl_C#G_0MsHo#RHRFVsl#_E0MsHo1Rrah)Qtz,Rh1) m pe7V_kH8GC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7kGVHC;89
R
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoR:aR1)tQh;RRRRRRRRRRRRRRRR-RR-HRLM$NsRs#0H
MoRRRR#CHx_#sCRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;RDRNHRN#VlsF_0L#soHMRRH#VlsF_s#0HRMor)1aQ,htR)zh p1me_ 7#GVHCR8
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0szMRh1) m pe7V_#H8GC9R;
RHNDNV#Rs_FlLNHMs#$_0MsHo#RHRFVsl0_#soHMRar1)tQh,hRz)m 1p7e _H#VG
C8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _H#VG9C8;R

RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRR:1Qa)hRt;RRRRRRRRRRRRRRRRRR--mNO0D0R#soHM
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
NRRD#HNRFVslO_F0_ND#H0sMHoR#sRVFFl_#H0sMroR1Qa)hRt,z h)1emp #7_VCHG8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp #7_VCHG8
9;
VRRk0MOHRFMVlsF_0E#soHMRR5
RERR#H0sMRoR:aR1)tQh;RRRRRRRRRRRRRRRR-RR-CREG0R#soHM
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
NRRD#HNRFVslC_EG0_#soHMRRH#VlsF_0E#soHMRar1)tQh,hRz)m 1p7e _H#VG
C8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp #7_VCHG8
9;
-RR-HR7s0CORMOFP#CsHRFMVOkM0MHF#R3R lGNb:DC
-RR-#RRHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-R-RkRV4<V=Rs_Fl#H0sM5oR"4j4jj34j;"2RR--n
36R-R-RRQM0#EHR#ONCER0C3R""#RHR0MFR0FbHNFMDN,RM08RE#CRHRxCFRV
RR--0RECFbk0kl0RkR#0lON0EGRCNDO0$R3
RR
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sM:oRR)1aQ2htRRRRRRRRRRRRRRRRR-RR-HRLM$NsRs#0H
MoRRRRskC0szMRh1) m pe7V_kH8GC;R
RNNDH#sRVFLl_#H0sMHoR#sRVF#l_0MsHo1Rrah)QtCRs0MksR)zh p1me_ 7kGVHC;89
NRRD#HNRFVslH_LM$Ns_s#0HRMoHV#Rs_Fl#H0sMroR1Qa)hstRCs0kMhRz)m 1p7e _HkVG9C8;R

RR--7CHsOF0ROD0NR8NMRGECRMOFP#CsHRFMVOkM0MHF#R3RQ0MRERH#OCN#
-RR-ER0C0R#soHMRMDCo#0ER#lk0NRl03OERGR NDlbCR:
RR--#MHoN#DRV:4R=VR#H8GCRR568MFI0-FRd
2;R-R-R4#VRR<=VlsF_0F#soHMR(5"4"3c2-R-R3-n6R
R
VRRk0MOHRFMVlsF_0F#soHMRR5
RFRR#H0sM:oRR)1aQ2htRRRRRRRRRRRRRRRRR-RR-ORm0RND#H0sMRo
RsRRCs0kMhRz)m 1p7e _HkVG;C8
NRRD#HNRFVslO_F0_ND#H0sMHoR#sRVFFl_#H0sMroR1Qa)hstRCs0kMhRz)m 1p7e _HkVG9C8;R

RMVkOF0HMsRVFEl_#H0sM5oR
RRRR0E#soHMR1:Rah)QtR2RRRRRRRRRRRRRRRRRRR--ERCG#H0sMRo
RsRRCs0kMhRz)m 1p7e _HkVG;C8
NRRD#HNRFVslC_EG0_#soHMRRH#VlsF_0E#soHMRar1)tQhR0sCkRsMz h)1emp k7_VCHG8
9;
VRRk0MOHRFMVlsF_s#0HRMo5R
RR#RL0MsHoRR:1Qa)hRt2RRRRRRRRRRRRRRRRR-R-RMLHNRs$#H0sMRo
RsRRCs0kMhRz)m 1p7e _H#VG;C8
NRRD#HNRFVsl#_L0MsHo#RHRFVsl0_#soHMRar1)tQhR0sCkRsMz h)1emp #7_VCHG8
9;RDRNHRN#VlsF_MLHN_s$#H0sMHoR#sRVF#l_0MsHo1Rrah)QtCRs0MksR)zh p1me_ 7#GVHC;89
R
RVOkM0MHFRFVsl#_F0MsHo
R5RRRRFs#0HRMo:aR1)tQh2RRRRRRRRRRRRRRRRRRR-m-ROD0NRs#0H
MoRRRRskC0szMRh1) m pe7V_#H8GC;R
RNNDH#sRVFFl_OD0N_s#0HRMoHV#Rs_FlFs#0HRMor)1aQRhtskC0szMRh1) m pe7V_#H8GC9
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHoRR:1Qa)hRt2RRRRRRRRRRRRRRRRR-R-RGECRs#0H
MoRRRRskC0szMRh1) m pe7V_#H8GC;R
RNNDH#sRVFEl_C#G_0MsHo#RHRFVsl#_E0MsHo1Rrah)QtCRs0MksR)zh p1me_ 7#GVHC;89
-
-RDs0_M#$0#ECHF#RM-
-RNbsoRlN#0$MEHC##M_F
M
C8NRbOo	NCHRVG_C8oCCMs_HOb;	o
H
DLssN$ RQ 
 ;kR#CQ   3avq] _)qNp3D
D;
ObN	CNoR8LF$HRVG_C8oCCMs_HObR	oHR#
RR--qEk0F7sRN8PHR#AHERFb5H8L#bEF@E@P8FD3s
o2R-R-REm0COsRFsM0H0LkC:s#RlKHRIpCHR#,YMNMHRO	toskMRH,)M$NRRW3]0HDFRM
RR--MDkDRsNsNO$RF0M#N#M0
ORRF0M#NRM0hwqzRz:Rh1) m pe7V_kH8GCRR5j8MFI04FR2=R:R05FE#CsRR=>'2j';R
RO#FM00NMR1hqwRR:z h)1emp #7_VCHG8jR5RI8FMR0F4:2R=FR50sEC#>R=R''j2R;
RMOF#M0N01Rhp:eRR71a_mzpt_QBea Bm5)RjFR8IFM0RR42:5=RFC0Es=#R>jR''
2;
-RR-ERaH8#RHCVVsRC8O#FM00NMRDIHDCR0D$DRFHkRVER0CNRbOo	NCFRL8H$R#$R#MC0E#NHxL
DCR-R-RRFsHDlbCMlC0RC8Ns#RCRNDMLklC,s#R0#CRR0F"k0sCH"RV$R#MC0E#NHxL3DC
ORRF0M#NRM0VCHG8M#$0FE_sC_sN:DRRmAmph qRR:=0Csk;R

RR--1ObCHRNDP#CsHRFMF"VRlHHMl"klRR0F8#FRFRlCLMFk8$NsRCOEOM	HoHRI0kEF0sRCs#Fs
VRRk0MOHRFMl#HMR,5DR:sRRaQh )t 2R
RRCRs0MksRaQh )t R
H#RCRLoRHMRR--VOkM0MHFRMlH#R
RRVRHRR5p=hRQa  t)F'DIsRFR=)RRaQh )t 'IDF2ER0CRM
RRRRR0sCkRsMjR;RRRRRRRRRRRRRRRRRRRRRR-RR-sRCsRFsO8FMHF0HM#,RHMDC0R
RRMRC8VRH;R
RRCRs0MksRMlHHllkR,5pR;)2
CRRMV8Rk0MOHRFMl#HM;R

RR--1ObCHRNDP#CsHRFMF"VRlHHMl"klRR0F8#FRFRlCLMFk8$NsRCOEOM	HoHRI0CERsssF#R
RVOkM0MHFRMlHCDR5,RRs:hRQa  t)R2
RsRRCs0kMhRQa  t)#RH
LRRCMoHR-R-RMVkOF0HMHRlMRC
RHRRVpR5RQ=Rhta  D)'FFIRsRR)=hRQa  t)F'DI02RE
CMRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&RRLzMF8kMCM8RkClLsNRb#8#C,NRI#RRNDCH0sRNDk8#C?R"
RRRRR#RRCsPCHR0$CFsssR;
RRRRR0sCkRsMjR;
RCRRMH8RVR;
RsRRCs0kMHRlMkHllpR5,2R);R
RCRM8VOkM0MHFRMlHC
;
R-R-RCaERDVFDHFIMVoRk0MOH#FMRCNsRCk#8MRFDH$RMs0CMDND$R3R sPC$kRVMHO0FRM
RR--ODND#OR"DMCNP"COR0CHERCs8CHsO$0DRRFsHHM8s0COD
$3R-R-RsbkbCF#:HRwGRC#"I8FM"0FRFbsLlDCR8NMR#sCFCDP#CRl0#NR0CN0#R
RVOkM0MHFRCODNCMPO
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-H-RM0bk
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)=R:RGlNHllk5oNs'VDC0N,Rsso'H0oE2R;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)=R:RMlH#s5NoC'DVR0,N'sosEHo0
2;RRRRPHNsNCLDR#sCkRD0RRRRRz:Rh1) m pe7V_#H8GCRs5NoN'sM2oC;R
RLHCoM-RR-kRVMHO0FOMRDMCNP
CORRRRNC##sM0RF50RN'soNC#OMM8HoMRN8NR5sDo'F/IR=hRQa  t)F'DI
22RRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRR&RRRe"RCFO0sNRb#8#CRHk#MNoRR0""FR""soNMCC,RGObC0RC8H"#R"I8FM"0F"R"
RRRRRP#CC0sH$sRCs;Fs
RRRR0sCkRsMN;so
CRRMV8Rk0MOHRFMONDCMOPC;R

RR--bbksF:#CRGwHC"#R8MFI0RF"bLsFDRClNRM8sFC#D#PCR0lCN0R#N#0C
VRRk0MOHRFMONDCMOPCRR5
RNRRs:oRR)zh p1me_ 7kGVHCR82RRRRRRRRR-RR-MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t RR:=lHNGl5klN'soD0CV,sRNoH'so2E0;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t RR:=l#HM5oNs'VDC0N,Rsso'H0oE2R;
RPRRNNsHLRDCskC#DR0RRRRR:hRz)m 1p7e _HkVGRC85oNs'MsNo;C2
LRRCMoHR-R-RMVkOF0HMDROCPNMCRO
RNRR#s#C0FRM0NR5sNo'#MOC8oHMR8NMRs5NoF'DI=R/RaQh )t 'IDF2R2
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRR&"CReOs0FR#bN#RC8kM#HoRRN"F"0"s"RNCMo,GRCb0COCH8R#"R"8MFI0"F""R
RRRRR#CCPs$H0RsCsF
s;RRRRskC0sNMRs
o;RMRC8kRVMHO0FOMRDMCNP;CO
R
R-a-R$RbCOPFMCRs0NkR"Mo#HM"C8R0HMFRRN"HkVG"C8,#RkCH8RMs0CMDND$R
RVOkM0MHFR_0FVCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7h_z1hQt R7;RR--#VEH0RC8P0COFRs
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)R;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RLHCoM-RR-kRVMHO0F0MRFH_VG
C8RRRRskC#D:0R=hRz)m 1p7e _HkVG5C8N2so;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0VF_H8GC;R

RR--aC$bRMOFP0CsR"NR#MHoCR8"HFM0RRNM"H#VG"C8,#RkCH8RMs0CMDND$R
RVOkM0MHFR_0FVCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;-RR-ER#HCV08CRPOs0F
RRRRMOF#M0N0CRDVH0_MG8CRRR:Q hat; )
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RCRLoRHMRR--VOkM0MHFR_0FVCHG8R
RRCRs#0kDRR:=z h)1emp #7_VCHG8s5No
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFR0_GVHC
8;
-RR-$RabOCRFCMPsN0RRV"kH8GC"MRH0NFRMkR"Mo#HM"C8,#RkCH8RMs0CMDND$R
RVOkM0MHFR_0FkRM#5R
RRsRNoRR:z h)1emp k7_VCHG8R2RRRRRRRRRR-R-RRVbP0COFRs
RsRRCs0kMhRz)m 1p7e _1zhQ th7R
RHR#
R#RRk$L0b0CRRRH#z h)1emp z7_ht1Qh5 7N'soEEHoRN-RsDo'F8IRF0IMF2Rj;R
RRNRPsLHND#CRD:PRR
0;RCRLoRHMRR--VOkM0MHFR_0Fk
M#RRRR#RDP:0=R5oNs2R;
RsRRCs0kMDR#PR;
R8CMRMVkOF0HMFR0_#kM;R

RR--aC$bRMOFP0CsRRNM"H#VG"C8R0HMFRRN"o#HM"C8,#RkCH8RMs0CMDND$R
RVOkM0MHFR_0F#
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-V-RbCRPOs0F
RRRR0sCkRsMz h)1emp 17_Q th7R
RHR#
R#RRk$L0b0CRRRH#z h)1emp 17_Q th7s5NoH'Eo-ERRoNs'IDFRI8FMR0Fj
2;RRRRPHNsNCLDRP#DR0:R;R
RLHCoM-RR-kRVMHO0F0MRF
_#RRRR#RDP:0=R5oNs2R;
RsRRCs0kMDR#PR;
R8CMRMVkOF0HMFR0_
#;
-RR-8RN84#RRR0F0RECpR1AF0VREMCRkClLsR
RbOsFCs8kCFRsk_M8k5bRNRsoRRRRRRR:HRMRz h)1emp k7_VCHG8R;
RRRRRRRRRRRRRRRRRRRRR#sCkRD0R:RRR0FkR)zh p1me_ 7kGVHC
8;RRRRRRRRRRRRRRRRRRRRRPRFCDsVFRIG:kRF0mRAmqp hH2R#R
RRNRPsLHNDNCRsMok#s,RCM#k#RR:z h)1emp z7_ht1QhR 75oNs'oEHEs-NoF'DIR+48MFI0jFR2R
RRRRR:5=RFC0Es=#R>jR''
2;RCRLoRHMRR--sMFk8b_k
RRRRoNskRM#5oNsk'M#EEHo-84RF0IMF2RjRR:=0kF_M5#RN2so;R
RRCRs##kMRRRRRRRRRRRRRRRRRRRRRRRRR=R:RoNskRM#+;R4
RRRR#sCkRD0:0=RFH_VG5C8skC#MN#5sEo'H-oEN'soD
FIRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFR8IFM0R,j2RoNs'oEHEN,RsDo'F;I2
RRRRCFPsFVDI:GR=sR5CM#k#C5s##kM'oEHE=2RR''42R;
R8CMRFbsOkC8ssCRF8kM_;kb
R
R-N-R8R8#4FR0RC0ERAp1RRFV0RECMLklCRs
RFbsOkC8ssCRF8kM_Rkb5oNsRRRRR:RRRRHMR)zh p1me_ 7#GVHC
8;RRRRRRRRRRRRRRRRRRRRRCRs#0kDRRRR:kRF0hRz)m 1p7e _H#VG;C8
RRRRRRRRRRRRRRRRRRRRFRRPVCsDGFIRF:RkA0Rm mpqRh2HR#
RPRRNNsHLRDCN#so,CRs#:#RR)zh p1me_ 71hQt 57RN'soEEHo-oNs'IDF+84RF0IMF2Rj;R
RLHCoM-RR-FRsk_M8kRb
RNRRsRo#5oNs#H'Eo4E-RI8FMR0Fj:2R=FR0_5#RN2so;R
RRsRNoN#5s'o#EEHo2RRRRRRRRRRRR=R:RoNs5oNs'oEHER2;RR--#MHoR0CGC
M8RRRRs#C#RRRRRRRRRRRRRRRRRRRRRRRR:N=RsRo#+;R4
RRRR#sCkRD0:0=RFH_VG5C8s#C#RC5s#E#'H-oE4R
RRRRRRRRRRRRRRRRRRRRRRRRRR8RRF0IMF2Rj,sRNoH'EoRE,N'soD2FI;R
RRPRFCDsVFRIG:5=R5oNs5oNs'oEHE/2R=CRs#s#5C'##EEHo-242
RRRRRRRRRRRRRRRRNRRM58RF5sR1_a7ztpmQeB_ mBa)C5s#2#2RR/='2j'2R;
R8CMRFbsOkC8ssCRF8kM_;kb
R
R-)-RF8kMHRMo-CRussVFlN#RRF"sk_M8MsCNC"#0R 5Q ( R6Rc2IOEHEFRsk#M8R
kbR-R-RCIEMER0CCRslMNH8RCsH>#RR6j33QRRVER0CCRslMNH8RCsQj1R306RERCMH0VRERC
RR--L0F0FLlRHH0R#RRN"R4"HH0R#FRskCM88F,R0sECICH#RRH0sNClHRM#0REC#CNl3R
RVOkM0MHFRksFMV8_H8GCRs5NoRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRRRRRRCRslMNH8RCsRRRRRz:Rh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDRksFMR8#RRRRRRRR:mRAmqp hR;
RPRRNNsHLRDCsMFk8P_FCDsVF:IRRmAmph q;R
RRNRPsLHNDsCRCD#k0RRRRRRRRRR:z h)1emp k7_VCHG8NR5sso'NCMo2R;
RoLCHRM
RsRRF8kM#=R:RDVN#
C;RRRRH5VRsNClHCM8sC'DMEo0R4>R2ER0CRM
RRRRRRHV5lsCN8HMC5sRsNClHCM8sH'EoRE2=4R''02RE
CMRRRRRRRRsMFk8:#R=NR5sNo5sDo'FRI2=4R''R2
RRRRRRRRRRRRRRRRRRFs5RFs5_0F#PkD5lsCN8HMCss5CHlNMs8C'oEHER-48MFI0RF
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRslMNH8'CsD2FI2=2RR''42R;
RRRRR8CMR;HV
RRRR#CDCR
RRRRRsMFk8:#R=NR5sNo5sDo'FRI2=4R''N2RM58RsNClHCM8ssR5CHlNMs8C'oEHE=2RR''42R;
RCRRMH8RVR;
RHRRVFRsk#M8RC0EMR
RRRRRsMFk8b_k5oNsRRRRR=RR>sRNoR,
RRRRRRRRRRRRRCRs#0kDRRRR=s>RCD#k0R,
RRRRRRRRRRRRRPRFCDsVFRIG=s>RF8kM_CFPsFVDI
2;RRRRCCD#
RRRRsRRCD#k0=R:RoNs;R
RRMRC8VRH;R
RRVRHRP5FCDsVF#I_0C$DRV=RH8GC_0#Nk0sNCN2RMs8RF8kM_CFPsFVDIER0CRM
RRRRR#sCkRD0:#=RNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRksFMV8_H8GC;R

RR--)MFk8oHMR#ONC0R#Nl0CC
M0RkRVMHO0FsMRF8kM_GVHC58RNRsoRRRRRRRRR:RRR)zh p1me_ 7#GVHC
8;RRRRRRRRRRRRRRRRRRRRRRRRsNClHCM8sRRRR:RRR)zh p1me_ 7#GVHC
8;RRRRRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRF8kM#RRRRRRRRRR:Apmm ;qh
RRRRsPNHDNLCFRsk_M8FsPCVIDFRA:Rm mpq
h;RRRRPHNsNCLDR#sCkRD0RRRRRRRR:hRz)m 1p7e _H#VGRC85oNs'MsNo;C2
LRRCMoH
RRRRksFMR8#:V=RNCD#;R
RRVRHRC5slMNH8'CsDoCM0>ERRR420MEC
RRRRHRRVsR5CHlNMs8CRC5slMNH8'CsEEHo2RR='24'RC0EMR
RRRRRRFRsk#M8RR:=5oNs5oNs'IDF2RR='24'
RRRRRRRRRRRRRRRRFRRsFR5s0R5Fk_#DsP5CHlNMs8C5lsCN8HMCEs'H-oE4FR8IFM0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsNClHCM8sF'DI222R'=R4;'2
RRRRCRRMH8RVR;
RCRRD
#CRRRRRFRsk#M8RR:=5oNs5oNs'IDF2RR='24'R8NMRC5slMNH8RCs5lsCN8HMCEs'H2oER'=R4;'2
RRRR8CMR;HV
RRRRRHVsMFk80#RE
CMRRRRRFRsk_M8kNb5sRoRRRRRRR=>N,so
RRRRRRRRRRRRRRRskC#DR0RR>R=R#sCk,D0
RRRRRRRRRRRRRRRFsPCVIDFG>R=RksFMF8_PVCsD2FI;R
RRDRC#RC
RRRRR#sCkRD0:N=Rs
o;RRRRCRM8H
V;RRRRHsVRF8kM_CFPsFVDIER0CRM
RRRRRRHV5CFPsFVDI0_#$RDC=HRVG_C8#kN0sCN02ER0CRM
RRRRRHRRVsRNos5NoH'EoRE2=jR''ER0CRM
RRRRRRRRR#sCkRD0:#=RNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;
RRRRRCRRD
#CRRRRRRRRRCRs#0kDRR:=MRF0#kN0sCN0RC5s#0kD'oEHEs,RCD#k0F'DI
2;RRRRRRRRCRM8H
V;RRRRRRRR-1-RHRoMLRH0MRF0VCHG8ERICIMRsbNbH
MoRRRRRMRC8VRH;R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMsMFk8H_VG;C8
R
R-O-RFCMPsR0#N#MRVCHG8MRH0NFRRHkVG3C8RERaCkRF00bkRRH#0REC#CNlRMDCoR0EN0#RERC
RR--HkMb0L,RCkON#NCRL"#54jjj"=2RRj"4jRj"=3RU
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRso:hRz)m 1p7e _H#VG2C8
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)=R:RoNs'oEHER;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)=R:RMlHCs5NoF'DIN,RsDo'F;I2
RRRRsPNHDNLCNRGsRoRRRRRRRR:z h)1emp #7_VCHG8C5DVH0_MG8C+84RF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDR#sCkRD0RRRRRz:Rh1) m pe7V_kH8GC5VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHVN'soDoCM0<ERR04RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RGRRNRsoR=R:R#NL5oNs2R;
RsRRCD#k0=R:R)zh p1me_ 7kGVHC58RGoNsRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FkGVHC
8;
------------------------------------------------------------------------------
-HRe#DHLCkRVMHO0F
M#-----------------------------------------------------------------------------R

RR--BPFMCHs#FVMRk0MOH#FM3aRRECC#RCNsRCMC8RC8VRFs#0$MEHC##ERICRsC0H$bODND$R
R-0-REFCRMRD$HkMb0MRN8kRF00bkRb0$C#RHR#NR0D8_FOoH_OPC03Fs
VRRk0MOHRFM0#F_kRDP5R
RRsRNoRR:z h)1emp k7_VCHG8R2RRRRRRRRRR-R-RGVHCb8RF0HMROPC0
FsRRRRskC0s1MRaz7_pQmtB _eB)am
HRR#R
RRNRPsLHNDsCRCD#k0RR:1_a7ztpmQeB_ mBa)NR5sDo'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVsRNoC'DMEo0R4<RRC0EMR
RRRRRskC0shMR1;pe
RRRR8CMR;HV
RRRR#sCkRD0:1=Raz7_pQmtB _eB)amRs5No
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFR0_D#kP
;
RkRVMHO0F0MRFk_#D5PR
RRRRoNsRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRRR--VCHG8FRbHRM0P0COFRs
RsRRCs0kMaR17p_zmBtQ_Be a
m)R#RH
RRRRsPNHDNLCCRs#0kDR1:Raz7_pQmtB _eB)amRs5NoC'DMEo0-84RF0IMF2Rj;R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR40MEC
RRRRsRRCs0kM1Rhp
e;RRRRCRM8H
V;RRRRskC#D:0R=aR17p_zmBtQ_Be aRm)5oNs2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0F#PkD;R

RMVkOF0HMFR0_P#DRR5
RNRRs:oRR)zh p1me_ 7kGVHCR82RRRRRRRRR-RR-HRVGRC8bMFH0CRPOs0F
RRRR0sCkRsM1_a7pQmtB _eB)amR
H#RCRLo
HMRRRRskC0s0MRFk_#DNP5s;o2
CRRMV8Rk0MOHRFM0#F_D
P;
VRRk0MOHRFM0#F_D5PR
RRRRoNsRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRRR--VCHG8FRbHRM0P0COFRs
RsRRCs0kMaR17m_pt_QBea BmH)R#R
RLHCoMR
RRCRs0MksR_0F#PkD5oNs2R;
R8CMRMVkOF0HMFR0_P#D;R

RMVkOF0HMFR0_HkVGRC85R
RRsRNoRRRRRRRRRRRRRRRR:RRR71a_mzpt_QBea BmR);RR--#VEH0RC8P0COFRs
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)R;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)R2
RsRRCs0kMMRksFC#D8PC_HkVG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RLHCoMR
RRVRHRs5NoC'DMEo0R4<RRRFssEHo0M_H8RCG>CRDVH0_MG8C2ER0CRM
RRRRR0sCkRsMhwqz;R
RRMRC8VRH;R
RRVRHRs5NoC'DMEo0RR/=skC#DD0'C0MoE02RE
CMRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNlR"&Razm_w QX7p51e"2R
RRRRRRRR"&Re0COFDsRC0MoE8#RFFRM0NRl03OERMRQbRk0DoCM0HER#
R"RRRRRRRR&hRQa  t)l'HN5oCN'soDoCM0RE2&RR"NRM8Fbk0kI0RHRDDL"CR
RRRRRRRRQ&Rhta  H)'lCNo5#sCk'D0DoCM0RE2&RR"ICH83R"
RRRRR#RRCsPCHR0$CFsssR;
RRRRR0sCkRsMhwqz;R
RRDRC#RC
RRRRR#sCkRD0:0=RFH_VGRC85oNsRRRRRRRRRR=>z h)1emp z7_ht1Qh5 7N2so,R
RRRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGR=D>RC_V0HCM8GR,
RRRRRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CRR=>sEHo0M_H82CG;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_HkVG;C8
R
RVOkM0MHFR_0F#GVHC58R
RRRRoNsRRRRRRRRRRRRRRRRRRR:1_a7ztpmQeB_ mBa)R;R-#-RE0HVCP8RCFO0sR
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t ;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t 2R
RRCRs0MksRskMCD#FP_C8#GVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5oNs'MDCoR0E<RR4FssRH0oE_8HMC>GRRVDC0M_H82CGRC0EMR
RRRRRskC0shMRq;1w
RRRR8CMR;HV
RRRRRHV5oNs'MDCoR0E/s=RCD#k0C'DMEo02ER0CRM
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_NRlC&aR"mw_1Q7X 5e1p2
R"RRRRRRRR&eR"CFO0sCRDMEo0#FR8R0MFR0lNORE3RbQMkD0RC0MoE#RHRR"
RRRRR&RRRaQh )t 'NHloNC5sDo'C0MoE&2RRN"RMF8Rkk0b0HRIDLDRC
R"RRRRRRRR&hRQa  t)l'HN5oCskC#DD0'C0MoE&2RRI"RH38C"R
RRRRRRCR#PHCs0C$RsssF;R
RRRRRskC0shMRq;1w
RRRR#CDCR
RRRRRskC#D:0R=FR0_GVHC58RNRsoRRRRRRRR=z>Rh1) m pe7Q_1t7h 5oNs2R,
RRRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRR=>D0CV_8HMC
G,RRRRRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8G>R=RosHEH0_MG8C2R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0F0MRFV_#H8GC;R

RR--a'IF#FROlCbDl0CMRlMkL,CsRFtsI0#REPCRCFO0s$RLRL4RH
03R-R-ROLCNCk#RL"N#4R5j3jjj2jjRj=R4jjj3jjj"sRFR#NL5n-42RR=4
n3RkRVMHO0F"MRN"L#RR5
RNRRs:oRR)zh p1me_ 7#GVHCR82RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t RR:=N'soEEHo;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t RR:=lCHM5oNs'IDF,sRNoF'DI
2;RRRRPHNsNCLDR#sC#RM#RRRRRz:Rh1) m pe7Q_1t7h Rs5NoC'DMEo0RI8FMR0Fj
2;RRRRPHNsNCLDR#sCkRD0RRRRRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8C+84RF0IMFHRso_E0HCM8G
2;RCRLo
HMRRRRH5VRN'soDoCM0<ERRF4RsCRs#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;1w
RRRR8CMR;HV
RRRR#sC#RM#5oNs'MDCo-0E4FR8IFM0RRj2:0=RFR_#5CODNCMPONR5s2o2;R
RRCRs###MRs5NoC'DMEo02RRRRRRRRRRRRR:=s#C#M5#RN'soDoCM04E-2R;R-C-RGMbN8HR#oLMRHR0
RsRRCD#k0RRRRRRRRRRRRRRRRRRRRRRRR=R:R_0FVCHG8NR5Ls#5CM###R2,D0CV_8HMC4G+,HRso_E0HCM8G
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMNR"L;#"
R
R-N-RDR#FoIsF#ER0CCRPOs0FRRL$4HRL0R3
RMVkOF0HM-R""
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)=R:RoNs'oEHE;+4
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hatR ):l=RH5MCN'soD,FIRoNs'IDF2R;
RPRRNNsHLRDCs#C#MR#RRRRR:hRz)m 1p7e _t1QhR 75oNs'MDCoR0E8MFI0jFR2R;
RPRRNNsHLRDCskC#DR0RRRRR:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5oNs'MDCoR0E<RR4FssRCD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRCRs###MRs5NoC'DMEo0-84RF0IMF2RjRR:=0#F_RD5OCPNMCNO5s2o2;R
RRCRs###MRs5NoC'DMEo02RRRRRRRRRRRRR:=s#C#M5#RN'soDoCM04E-2R;R-C-RGMbN8HR#oLMRHR0
RsRRCD#k0RRRRRRRRRRRRRRRRRRRRRRRR=R:R_0FVCHG8-R5s#C#MR#,D0CV_8HMCRG,sEHo0M_H82CG;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM";-"
R
R-q-R808HH
FMRkRVMHO0F"MR+5"R
RRRRRD,sRR:z h)1emp k7_VCHG8R2RR-R-RHkVG5C8NFR8IFM0RRL2+VRkH8GC58ORF0IMF2R8RR=
RsRRCs0kMhRz)m 1p7e _HkVGRC8RRRR-k-RVCHG8N5lG,5NO42+RI8FMR0Fl5HML2,82R
RHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2;+4
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=lCHM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCskC#DR0RRRRRRRRRRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRR:z h)1emp z7_ht1QhR 75VDC0M_H8-CGsEHo0M_H8
CGRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0D_#PRR:z h)1emp z7_ht1QhR 75VDC0M_H8-CGsEHo0M_H8
CGRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRF0IMF2Rj;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRF4RsCRs#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;zw
RRRR8CMR;HV
RRRRCDs#CHxRRRR:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxCR:RR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RDRR#RDPRRRRR=R:R_0FkRM#5CDs#CHx2R;
RsRR#RDPRRRRR=R:R_0FkRM#5Css#CHx2R;
RsRRCD#k0D_#P=R:RDD#PRR+sP#D;R
RRCRs#0kDRRRRRR:=0VF_H8GC5#sCk_D0#,DPRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR""+;R

RMVkOF0HM+R""
R5RRRRDs,RRz:Rh1) m pe7V_#H8GC2RRRRR--#GVHCN85RI8FMR0FL+2RRH#VG5C8OFR8IFM0RR82=RR
RsRRCs0kMhRz)m 1p7e _H#VGRC8RRRR-#-RVCHG8N5lG,5NO42+RI8FMR0Fl5HML2,82R
RHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2;+4
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=lCHM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp #7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCskC#DR0RRRRRRRRRRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _t1QhR 75VDC0M_H8-CGsEHo0M_H8RCG8MFI0jFR2R;
RPRRNNsHLRDCskC#D#0_DRPRRRRRRz:Rh1) m pe7Q_1t7h RC5DVH0_MG8C-osHEH0_MG8CRI8FMR0Fj
2;RCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<RRRFsskC#DD0'C0MoERR<402RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RDRRsHC#xRCRR=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HCRRRRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDD#PRRRRRRR:0=RFR_#5CDs#CHx2R;
RsRR#RDPRRRRR=R:R_0F#sR5sHC#x;C2
RRRR#sCk_D0#RDP:D=R#RDP+#RsD
P;RRRRskC#DR0RR:RR=FR0_GVHCs85CD#k0D_#PD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MR+
";
-RR-kR1LN0sOF0HMR
RVOkM0MHFR""-RR5
RDRR,RRs:hRz)m 1p7e _HkVG2C8RRRR-k-RVCHG8R5N8MFI0LFR2RR-kGVHCO85RI8FMR0F8=2R
RRRR0sCkRsMz h)1emp k7_VCHG8RRRR-R-RHkVG5C8l5NGN2,O+84RF0IMFHRlM,5L8
22R#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo+E24R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMDC5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLCCRs#0kDRRRRRRRRR:RRR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDP:hRz)m 1p7e _1zhQ th7DR5C_V0HCM8GH-so_E0HCM8GR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2;RRRRPHNsNCLDR#sCk_D0#RDP:hRz)m 1p7e _1zhQ th7DR5C_V0HCM8GH-so_E0HCM8GR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2;RCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<RRRFsskC#DD0'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RDRRsHC#xRCRR=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HCRRRRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDD#PRRRRRRR:0=RFM_k#DR5sHC#x;C2
RRRRDs#PRRRRRRR:0=RFM_k#sR5sHC#x;C2
RRRR#sCk_D0#RDP:D=R#RDP-#RsD
P;RRRRskC#DR0RR:RR=FR0_GVHCs85CD#k0D_#PD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MR-
";
VRRk0MOHRFM"R-"5R
RR,RDR:sRR)zh p1me_ 7#GVHCR82R-RR-VR#H8GC58NRF0IMF2RLR#-RVCHG8R5O8MFI08FR2RR=
RRRR0sCkRsMz h)1emp #7_VCHG8RRRR-R-RH#VG5C8l5NGN2,O+84RF0IMFHRlM,5L8
22R#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo+E24R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMDC5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLCCRs#0kDRRRRRRRRR:RRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5C_V0HCM8GH-so_E0HCM8GFR8IFM0R;j2
RRRRsPNHDNLCCRs#0kD_P#DRRRRR:RRR)zh p1me_ 71hQt 57RD0CV_8HMCsG-H0oE_8HMC8GRF0IMF2Rj;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRF4RsCRs#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;1w
RRRR8CMR;HV
RRRRCDs#CHxRRRR:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxCR:RR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RDRR#RDPRRRRR=R:R_0F#DR5sHC#x;C2
RRRRDs#PRRRRRRR:0=RFR_#5Css#CHx2R;
RsRRCD#k0D_#P=R:RDD#PRR-sP#D;R
RRCRs#0kDRRRRRR:=0VF_H8GC5#sCk_D0#,DPRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR""-;R

RMVkOF0HM*R""
R5RRRRDs,RRz:Rh1) m pe7V_kH8GC2RRRRR--kGVHCN85RI8FMR0FL*2RRHkVG5C8OFR8IFM0RR82=R
RRCRs0MksR)zh p1me_ 7kGVHCR8RR-RR-VRkH8GC5ON++84RF0IMF+RL8R2
R
H#RRRRPHNsNCLDRDD#PRRRRRRR:hRz)m 1p7e _1zhQ th7DR5'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLC#RsDRPRRRRRRz:Rh1) m pe7h_z1hQt 57RsC'DMEo0-84RF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0D_#PRR:z h)1emp z7_ht1QhR 75Ds'C0MoE'+DDoCM04E-RI8FMR0Fj
2;RRRRPHNsNCLDR#sCkRD0RRRR:hRz)m 1p7e _HkVGRC85ED'HRoE+'RsEEHo+84RF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlRRH5MCDF'DID,R'IDF2RR+lCHM5Ds'FRI,sF'DI;22
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<4sRF
RRRRRRRR#sCk'D0DoCM0/ER=CRs#0kD_P#D'MDCo20ERC0EMR
RRRRRskC0shMRq;zw
RRRR8CMR;HV
RRRRDD#PRRRRRRR:0=RFM_k#OR5DMCNP5COD;22
RRRRDs#PRRRRRRR:0=RFM_k#OR5DMCNP5COs;22
RRRR#sCk_D0#RDP:D=R#RDP*#RsD
P;RRRRskC#DR0RR:RR=FR0_GVHC58RskC#D#0_DRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM";*"
R
RVOkM0MHFR""*RR5
RDRR,RRs:hRz)m 1p7e _H#VG2C8RRRR-#-RVCHG8R5N8MFI0LFR2RR*#GVHCO85RI8FMR0F8=2RRR
RRCRs0MksR)zh p1me_ 7#GVHCR8RR-RR-VR#H8GC5ON++84RF0IMF+RL8R2
R
H#RRRRPHNsNCLDRDD#PRRRRRRR:hRz)m 1p7e _t1QhR 75DD'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCsP#DRRRRR:RRR)zh p1me_ 71hQt 57RsC'DMEo0-84RF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0D_#PRR:z h)1emp 17_Q th7sR5'MDCo+0EDC'DMEo0-84RF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0RRRRRR:z h)1emp #7_VCHG8DR5'oEHERR+sH'Eo4E+RI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMlHC'5DD,FIRDD'FRI2+HRlMsC5'IDF,'RsD2FI2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<RR4FRs
RRRRRsRRCD#k0C'DMEo0RR/=skC#D#0_DDP'C0MoE02RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RDRR#RDPRRRRR=R:R_0F#OR5DMCNP5COD;22
RRRRDs#PRRRRRRR:0=RFR_#5CODNCMPO25s2R;
RsRRCD#k0D_#P=R:RDD#PRR*sP#D;R
RRCRs#0kDRRRRRR:=0VF_H8GCRC5s#0kD_P#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HM*R""
;
RkRVMHO0F"MR/5"R
RRRRRD,sRR:z h)1emp k7_VCHG8R2RR-R-RHkVG5C8NFR8IFM0RRL2/VRkH8GC58ORF0IMF2R8R
=RRRRRskC0szMRh1) m pe7V_kH8GCRRH#RRRRRRRR-R-RkGVHCN85-88RF0IMF-RLO2-4
LRRCMoH
RRRR0sCkRsM8HHP85CRDs,R2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MR/5"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RR-R-RH#VG5C8NFR8IFM0RRL2/VR#H8GC58ORF0IMF2R8R
=RRRRRskC0szMRh1) m pe7V_#H8GCRRH#RRRRRRRR-#-RVCHG8-5N8R+48MFI0LFR-
O2RCRLo
HMRRRRskC0s8MRH8PHCDR5,2Rs;R
RCRM8VOkM0MHFR""/;R

RR--a#EHRsPC#MHFRRFV8HHP8oCRH#PCRC0ERCk#sFRlsOCRFsM0FRD
RR--kGVHCN85RI8FMR0FL/2RRHkVG5C8OFR8IFM0RR82=VRkH8GC58N-RI8FMR0FL--O4R2
RMVkOF0HMHR8PCH8RR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8
RRRRMOF#M0N0FRsk_M8#D0$CRR:VCHG8F_sk_M8#D0$C$_0b:CR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRR:hzqa)RqpRRRRRRRRRRRRR:RR=HRVG_C8oskN8H_L0
#2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDsCRCD#k0RRRRRR:z h)1emp k7_VCHG8DR5'oEHERR-lCHM5Ds'FRI,sF'DI82RF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlRRHRMC5DD'FRI,DF'DI-2RREs'HRoE-;42
RRRRsPNHDNLCsR8CD#k0RRRRz:Rh1) m pe7V_kH8GCRC5s#0kD'oEHEFR8IFM0R#sCk'D0DRFI-NoksL8_H20#;R
RRNRPsLHNDDCRsHC#xRCRRRR:z h)1emp k7_VCHG8DR5'oEHEFR8IFM0RED'HRoE-sR8CD#k0C'DMEo0+;42
RRRRsPNHDNLC#RDDRPRRRRRRz:Rh1) m pe7h_z1hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RRRRPHNsNCLDRDs#PRRRRRRR:hRz)m 1p7e _1zhQ th7sR5'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kD_P#DRz:Rh1) m pe7h_z1hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<RR
FsRRRRRRRRl#HM5Ds'FRI,sF'DI/2R='RsDRFIFlsRH5M#DF'DID,R'IDF2=R/RDD'FRI20MEC
RRRRsRRCs0kMqRhz
w;RRRRCRM8H
V;RRRRD#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R
D,RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=RCDs#CHx'oEHER,
RRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>D#sCH'xCD,FI
RRRRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D=CR>HRVG_C8IbsN,RRR-P-RCFO0sMRFDo$Rs#FI
RRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>HRVG_C80MskOCN02R;
RDRR#RDP:0=RFM_k#OR5DMCNPRCO5CDs#CHx2
2;RRRRsP#DRR:=0kF_M5#RONDCMOPCR25s2R;
RHRRVsR5#RDP=2RjRC0EMR
RRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRRQ"7e Q75HkVG2C8RP7HHF#HM$RLRsxCF#"RCsPCHR0$CFsssR;
RRRRR#sCkRD0:#=RNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;RR-R-R0#Nk0sNCR
RRDRC#RC
RRRRR#sCk_D0#RDP:D=R#RDP/#RsD
P;RRRRRsR8CD#k0RRRRR:=0VF_H8GCRC5s#0kD_P#D,sR8CD#k0H'EoRE,8#sCk'D0D2FI;R
RRRRRskC#D:0R=CRs#CHxRs5NoRRRRRRRRRRRRR=>8#sCk,D0
RRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=s>RCD#k0H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>CRs#0kD'IDF,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>VCHG8s_INRb,RR--FsPCVIDFRbHlFH##L
DCRRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$C
2;RRRRCRM8H
V;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMHR8PCH8;R

RR--#GVHCN85RI8FMR0FL/2RRH#VG5C8OFR8IFM0RR82=VR#H8GC58N-+84RF0IMF-RLOR2
RMVkOF0HMHR8PCH8RR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8
RRRRMOF#M0N0FRsk_M8#D0$CRR:VCHG8F_sk_M8#D0$C$_0b:CR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRR:hzqa)RqpRRRRRRRRRRRRR:RR=HRVG_C8oskN8H_L0
#2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RRRRRR:z h)1emp #7_VCHG8DR5'oEHERR-lCHM5Ds'FRI,sF'DI+2RR84RF0IMFRR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlCHMR'5DD,FIRDD'FRI2-'RsEEHo2R;
RPRRNNsHLRDC8#sCkRD0R:RRR)zh p1me_ 7#GVHC58RskC#DE0'HRoE8MFI0sFRCD#k0F'DIk-oN_s8L#H02R;
RPRRNNsHLRDCD#sCHRxCR:RRR)zh p1me_ 7#GVHC58RDH'Eo4E+RI8FMR0FDH'Eo4E+Rs-8CD#k0C'DMEo0+;42
RRRRsPNHDNLC#RDDRPRRRRRRz:Rh1) m pe7Q_1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RRNRPsLHNDsCR#RDPRRRRRRR:z h)1emp 17_Q th7sR5'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kD_P#DRz:Rh1) m pe7Q_1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRF4RsR
RRRRRRHRlMs#5'IDF,'RsD2FIRR/=sF'DIsRFRMlH#'5DD,FIRDD'FRI2/D=R'IDF2ER0CRM
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=D>R,R
RRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=D>RsHC#xEC'H,oE
RRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>sRDCx#HCF'DIR,
RRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>VCHG8s_INRb,R-R-ROPC0RFsF$MDRFosIR#
RRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>VCHG8s_0kNMO0;C2
RRRRDD#P=R:R_0F#OR5DMCNPRCO5CDs#CHx2
2;RRRRsP#DRR:=0#F_RD5OCPNMC5ORs;22
RRRRRHV5Ds#PRR=j02RE
CMRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R7QQe7# 5VCHG872RH#PHHRFMLx$RC"sFRP#CC0sH$sRCs;Fs
RRRRsRRCD#k0=R:R0#Nk0sNCsR5CD#k0H'EoRE,skC#DD0'F;I2
RRRR#CDCR
RRRRRskC#D#0_D:PR=#RDD/PRRDs#PR;
RRRRRC8s#0kDRRRR:0=RFH_VGRC85#sCk_D0#,DPRC8s#0kD'oEHE8,RskC#DD0'F;I2
RRRRsRRCD#k0=R:R#sCHRxC5oNsRRRRRRRRRRRR=8>RskC#D
0,RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>CRs#0kD'oEHER,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=R#sCk'D0D,FI
RRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=V>RH8GC_NIsbR,R-F-RPVCsDRFIHFlb#L#HDRC
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D2R;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRP8HH;8C
R
R-4-RRk/RVCHG8R5N8MFI0LFR2RR=kGVHC-85LFR8IFM0R--N4R2
RMVkOF0HMCRsOsHbFDONRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMRCFMRz:Rh1) m pe7V_kH8GCRR5j8MFI0jFR2=R:R""4;R
RLHCoMR
RRCRs0MksRP8HHR8C5RDRRRRRRRRRRR=>F,MC
RRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRkRoN_s8L#H0R>R=RNoksL8_H20#;R
RCRM8VOkM0MHFROsCHFbsO;ND
R
R-4-RR#/RVCHG8R5N8MFI0LFR2RR=#GVHC-85LR+48MFI0-FRNR2
RMVkOF0HMCRsOsHbFDONRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRO#FM00NMRCFMRRRRRz:Rh1) m pe7V_#H8GCRR548MFI0jFR2=R:R4"j"R;R-C-RGN0sR0LH3R
RRNRPsLHNDsCRCD#k0:GRR)zh p1me_ 7#GVHC58R-MlHCs5NoF'DIN,RsDo'F+I2.FR8IFM0Rs-NoH'Eo;E2
LRRCMoH
RRRRRHV5oNs'MDCoR0E<RR4FssRCD#k0DG'C0MoERR<402RE
CMRRRRRCRs0MksR1hqwR;
RCRRD
#CRRRRRCRs#0kDG=R:RP8HHR8C5RDRRRRRRRRRRR=>F,MC
RRRRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRoskN8H_L0R#R=o>Rk8Ns_0LH#
2;RRRRRCRs0MksR#sCkGD0RC5s#0kDGH'Eo4E-RI8FMR0FskC#D'0GD2FI;-RR-CRslCFPR0CGsLNRHR0
RCRRMH8RVR;
R8CMRMVkOF0HMCRsOsHbFDON;R

RR--kGVHC58RNFR8IFM0RRL2sRClkGVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VRkH8GCRH5lM,5NO82RF0IMFHRlM,5L8
22RkRVMHO0F"MRs"ClRR5
RDRR,RRs:hRz)m 1p7e _HkVG2C8RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0ssMRCHlNMs8CR,5DR;s2
CRRMV8Rk0MOHRFM"lsC"
;
R-R-RlsCN8HMCRs
RR--#GVHC58RNFR8IFM0RRL2sRCl#GVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VR#H8GCRH5lM,5NO82RF0IMFHRlM,5L8
22RkRVMHO0F"MRs"ClRR5
RDRR,RRs:hRz)m 1p7e _H#VG2C8RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0ssMRCHlNMs8CR,5DR;s2
CRRMV8Rk0MOHRFM"lsC"
;
R-R-RHkVGRC858NRF0IMF2RLRlsCRHkVGRC858ORF0IMF2R8
-RR-RRRRRRRRk=RVCHG8lR5HNM5,RO28MFI0lFRHLM5,282
VRRk0MOHRFMsNClHCM8s
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRFROMN#0Ms0RF8kM_$#0D:CRRGVHCs8_F8kM_$#0D0C_$RbC:V=RH8GC_ksFM#8_0C$D;R
RRFROMN#0Mo0Rk8Ns_0LH#:RRRahqzp)qRRRRRRRRRRRRRRRR:V=RH8GC_NoksL8_H20#
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RPRRNNsHLRDCskC#DR0RR:RRR)zh p1me_ 7kGVHC58RlHHMl5klDH'EoRE,sH'EoRE28MFI0RF
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlCHM5DD'FRI,sF'DI;22
RRRRsPNHDNLCsRDCx#HCRRRRz:Rh1) m pe7V_kH8GCRN5lGkHll'5DEEHo,'RsD2FIRI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMlH#'5sD,FIRDs'F-I2oskN8H_L0;#2
RRRRsPNHDNLCsRsCx#HCRRRRz:Rh1) m pe7V_kH8GCR'5sEEHoRI8FMR0FsF'DIk-oN_s8L#H02R;
RPRRNNsHLRDC8#sCkRD0R:RRR)zh p1me_ 7kGVHC58Rs#sCH'xCsoNMC
2;RRRRPHNsNCLDRDD#PRRRRRRR:hRz)m 1p7e _1zhQ th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCsP#DRRRRR:RRR)zh p1me_ 7zQh1t7h Rs5sCx#HCC'DMEo0-84RF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0D_#PRR:z h)1emp z7_ht1QhR 75Ds#PN'sM2oC;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRF4RsR
RRRRRRHRlMs#5'IDF,'RsD2FIRR/=sF'DIsRFRMlH#'5DD,FIRDD'FRI2/D=R'IDF2ER0CRM
RRRRR0sCkRsMhwqz;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=D>R,R
RRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=D>RsHC#xEC'H,oE
RRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>sRDCx#HCF'DIR,
RRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>VCHG8s_INRb,RRRR-P-RCFO0sMRFDo$Rs#FI
RRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>HRVG_C80MskOCN02R;
RDRR#RDP:0=RFM_k#DR5sHC#x;C2
RRRRCss#CHxRR:=sHC#x5CRNRsoRRRRRRRRR=RR>,Rs
RRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>sRsCx#HCH'Eo
E,RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=RCss#CHx'IDF,R
RRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=V>RH8GC_NIsbR,RR-RR-CRPOs0FRDFM$sRoF
I#RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RGVHC08_sOkMN20C;R
RR#RsD:PR=FR0_#kMRs5sCx#HC
2;RRRRH5VRsP#DRj=R2ER0CRM
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&sR"CHlNMs8C5HkVG2C8RP7HHF#HM$RLRsxCF#"RCsPCHR0$CFsssR;
RRRRR#sCkRD0:#=RNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;RRRRR-#-RNs0kN
0CRRRRCCD#
RRRRHRRVsR5'IDFRR<=DH'EoRE20MEC
RRRRRRRR#sCk_D0#RDP:D=R#RDPsRClsP#D;R
RRRRRRsR8CD#k0RRRRR:=0VF_H8GCRC5s#0kD_P#D,sR8CD#k0H'EoRE,8#sCk'D0D2FI;R
RRRRRRCRs#0kDRR:=sHC#x5CRNRsoRRRRRRRRR=RR>sR8CD#k0R,
RRRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=s>RCD#k0H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>skC#DD0'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>VCHG8s_INRb,RR--O'NM0PRFCDsVFRI
RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D;C2
RRRRCRRMH8RVR;
RRRRRRHVDF'DIRR<sF'DIER0CRM
RRRRRsRRCD#k0H5lMs#5'IDF-R4,DH'EoRE28MFI0DFR'IDF2=R:
RRRRRRRRORRDMCNP5CODH5lMs#5'IDF-R4,DH'EoRE28MFI0DFR'IDF2
2;RRRRRMRC8VRH;R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMsNClHCM8s
;
R-R-RlsCN8HMCRs
RR--#GVHC58RNFR8IFM0RRL2sRCl#GVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VR#H8GCRH5lM,5NO82RF0IMFHRlM,5L8
22RkRVMHO0FsMRCHlNMs8CRR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RGVHCb8RF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:HRVG_C8sMFk80_#$_DC0C$bRR:=VCHG8F_sk_M8#D0$CR;
RORRF0M#NRM0oskN8H_L0R#R:qRhaqz)pRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRPHNsNCLDRND_LR#RRRRR:hRz)m 1p7e _HkVGRC85sD'NCMo2R;
RPRRNNsHLRDCsL_N#RRRR:RRR)zh p1me_ 7kGVHC58RsN'sM2oC;R
RRNRPsLHNDsCRCD#k0RRRRRR:z h)1emp #7_VCHG8lR5HlMHksl5'oEHED,R'oEHE82RF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlRRH5MCsF'DID,R'IDF2
2;RRRRPHNsNCLDRoMC_#sCkRD0:hRz)m 1p7e _H#VGRC85MlHHllk5Es'H,oERED'H2oE+84RF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlRRH5M#sF'DID,R'IDF2
2;RCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<RR
FsRRRRRRRRl#HM5Ds'FRI,sF'DI/2R='RsDRFIFlsRH5M#DF'DID,R'IDF2=R/RDD'FRI20MEC
RRRRsRRCs0kMqRh1
w;RRRRCRM8H
V;RRRRDL_N#=R:R_0FkGVHC58RD
2;RRRRsL_N#=R:R_0FkGVHC58Rs
2;RRRRskC#D:0R=hRz)m 1p7e _H#VGRC85lsCN8HMC5sR
RRRRDRRRRRRRRRRR=RR>_RDN,L#
RRRRsRRRRRRRRRRR=RR>_RsN,L#
RRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$C;22
RRRRoMC_#sCkRD0:-=RskC#D
0;RRRRHDVR5ED'H2oER'=R40'RE
CMRRRRRCRs#0kDRR:=M_CoskC#Ds05CD#k0N'sM2oC;R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMsNClHCM8s
;
R-R-R8lFk
DFR-R-RHkVGRC858NRF0IMF2RLR8lFRHkVGRC858ORF0IMF2R8
-RR-RRRRRRRRk=RVCHG8lR5HNM5,RO28MFI0lFRHLM5,2R82R
RVOkM0MHFRF"l85"R
RRRRRD,sRR:z h)1emp k7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksR8lFkRDF5RD,s
2;RMRC8kRVMHO0F"MRl"F8;R

RR--#GVHC58RNFR8IFM0RRL2lRF8#GVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VR#H8GCRR5O8MFI0lFRHLM5,2R82R
RVOkM0MHFRF"l85"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksR8lFk5DFDs,R2R;
R8CMRMVkOF0HMlR"F;8"
R
R-l-RFD8kFR
R-k-RVCHG8NR5RI8FMR0FLl2RFk8RVCHG8OR5RI8FMR0F8R2
RR--RRRRR=RRRHkVGRC85MlH5ON,2FR8IFM0RMlH5RL,8
22RkRVMHO0FlMRFD8kF
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRV:RH8GC_ksFM#8_0C$D_b0$C=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#Rh:Rq)azqRpRRRRRRRRRRRRRR=R:RGVHCo8_k8Ns_0LH#R2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMCRslMNH85CsDRRRRRRRRRRR=D>R,R
RRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=RR>,Rs
RRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$C>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRoRRk8Ns_0LH#=RR>kRoN_s8L#H02R;
R8CMRMVkOF0HMFRl8FkD;R

RR--#GVHC58RNFR8IFM0RRL2lRF8#GVHC58ROFR8IFM0R
82R-R-RRRRRRRR=VR#H8GCRR5O8MFI0lFRHLM5,2R82R
RVOkM0MHFR8lFkRDF5R
RR,RDRRsRRRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-V-RH8GCRHbFMH0RM0bk
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#RRRR:qRhaqz)pRRRRRRRRRRRRRRRRRRR:V=RH8GC_NoksL8_H20#
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCDL_N#RR:z h)1emp k7_VCHG8DR5'MsNo;C2
RRRRsPNHDNLC_RsNRL#:hRz)m 1p7e _HkVGRC85ss'NCMo2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RsH'Eo8ERF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlRRH5MCsF'DID,R'IDF2
2;RRRRPHNsNCLDRC8s#0kDRz:Rh1) m pe7V_#H8GCRH5lMkHll'5sEEHo,'RDEEHo2R+48MFI0RF
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMlH#'5sD,FIRDD'F2I2;R
RRNRPsLHND8CRskC#DM0_Fx0_CRsF:mRAmqp hR;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<RR4FRs
RRRRRlRRH5M#sF'DIs,R'IDF2=R/RDs'FFIRsHRlMD#5'IDF,'RDD2FIRR/=DF'DI02RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RDRR_#NLRR:=0kF_VCHG8DR52R;
RsRR_#NLRR:=0kF_VCHG8sR52R;
R8RRskC#D:0R=jR""RR&z h)1emp #7_VCHG8C5slMNH8RCs5RDRRRRRRRRRRR=>DL_N#R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=>sL_N#R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRR=>sMFk80_#$2DC2R;
RHRRV0R5F5_#8#sCk2D0Rj=R2ER0CRM
RRRRRC8s#0kD_0MF_sxCF=R:RDVN#
C;RRRRCCD#
RRRR8RRskC#DM0_Fx0_CRsF:0=Rs;kC
RRRR8CMR;HV
RRRRRHV0GF_jD455ED'H2oE2RR='R4'NRM80GF_js455Es'H2oE2RR='
j'RRRRRMRN8sR8CD#k0F_M0C_xs0FRE
CMRRRRRCRs#0kDRR:=sHC#x5CRNRsoRRRRRRRRR=RR>RRs-sR8CD#k0R,
RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=R#sCk'D0EEHo,R
RRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>skC#DD0'F
I,RRRRRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D=CR>PRFCDsVF#I_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$2DC;R
RRDRC#RHV0GF_jD455ED'H2oE2RR='R4'NRM80GF_js455Es'H2oE2RR='R4'0MEC
RRRRsRRCD#k0=R:R#sCHRxC5oNsRRRRRRRRRRRR=->R8#sCk,D0
RRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=s>RCD#k0H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>CRs#0kD'IDF,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$C
2;RRRRCHD#VFR0_4Gj5DD5'oEHER22=jR''MRN8FR0_4Gj5ss5'oEHER22=4R''R
RRRRRNRM88#sCk_D0M_F0xFCsRC0EMR
RRRRRskC#D:0R=CRs#CHxRs5NoRRRRRRRRRRRRR=>8#sCkRD0+,Rs
RRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=s>RCD#k0H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>CRs#0kD'IDF,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$C
2;RRRRCCD#
RRRRsRRCD#k0=R:R#sCHRxC5oNsRRRRRRRRRRRR=8>RskC#D
0,RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>CRs#0kD'oEHER,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=R#sCk'D0D,FI
RRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$CR,
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D2R;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR8lFk;DF
R
R-u-RsCFO8CksRsVFRF0E#ICREMFRCRC8N"MRNkOOlNkD0"FsRMVkOF0HMR
RbOsFCs8kC8RN8N_OsRs$5R
RR,RpRR)RRH:RMzRRh1) m pe7V_kH8GC;R
RR_ROHRMRRH:RM1RRaz7_pQmtBR;
RsRRCD#k0RR:FRk0z h)1emp k7_VCHG8R;
RORR_0FkRRR:FRk01_a7ztpmQRB2HR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2;+4
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=l#HM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCDP#D,#RsD:PRR)zh p1me_ 7zQh1t7h RC5DVH0_MG8C-osHEH0_MG8C
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2R;
RPRRNNsHLRDCskC#D#0_D:PRR)zh p1me_ 7zQh1t7h RC5DVH0_MG8C-osHEH0_MG8C
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2R;
RPRRNNsHLRDCO:GRR)zh p1me_ 7zQh1t7h RR5j8MFI0jFR2R;R-B-RN$ssR
HMRCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<R2ER0CRM
RRRRR#sCkRD0:h=Rq;zw
RRRRORR_0FkR=R:R''j;R
RRDRC#RC
RRRRRROG5Rj2RRRR:O=R_;HM
RRRRDRRsHC#xRCRR=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRs#sCHRxCR:RR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRRRR:0=RFM_k#DR5sHC#x;C2
RRRRsRR#RDPRRRRR=R:R_0FkRM#5Css#CHx2R;
RRRRR#sCk_D0#RDP:D=R#RDP+#RsD+PRR;OG
RRRRORR_0FkRRRRR=R:R#sCk_D0#5DPD0CV_8HMC;G2
RRRRsRRCD#k0=R:R_0FVCHG8C5s#0kD_P#DRC5DVH0_MG8C-osHEH0_MG8C-84RF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8G,-4RosHEH0_MG8C2R;
RCRRMH8RVR;
R8CMRFbsOkC8sNCR8O8_N$ss;R

RFbsOkC8sNCR8O8_N$ssRR5
RpRR,RR)RRR:HRMRz h)1emp #7_VCHG8R;
RORR_RHMRRR:HRMR1_a7ztpmQ
B;RRRRskC#D:0RR0FkR)zh p1me_ 7#GVHC
8;RRRROk_F0:RRR0FkR71a_mzpt2QBR
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE42+;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDP:hRz)m 1p7e _t1QhR 75VDC0M_H8-CGsEHo0M_H8
CGRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2;RRRRPHNsNCLDR#sCk_D0#RDP:hRz)m 1p7e _t1QhR 75VDC0M_H8-CGsEHo0M_H8
CGRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2;RRRRPHNsNCLDRROG:hRz)m 1p7e _t1QhR 7584RF0IMF2Rj;-RR-NRBsRs$HRM
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRskC#D:0R=qRh1
w;RRRRR_ROFRk0RR:=';j'
RRRR#CDCR
RRRRRO5GR4R2RR:RR=jR''R;
RRRRRROG5Rj2RRRR:O=R_;HM
RRRRDRRsHC#xRCRR=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRs#sCHRxCR:RR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRRRR:0=RFR_#5CDs#CHx2R;
RRRRRDs#PRRRRRRR:0=RFR_#5Css#CHx2R;
RRRRR#sCk_D0#RDP:D=R#RDP+#RsD+PRR;OG
RRRRORR_0FkRRRRR=R:R#sCk_D0#5DPD0CV_8HMC;G2
RRRRsRRCD#k0=R:R_0FVCHG8C5s#0kD_P#DRC5DVH0_MG8C-osHEH0_MG8C-84RF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8G,-4RosHEH0_MG8C2R;
RCRRMH8RVR;
R8CMRFbsOkC8sNCR8O8_N$ss;R

RR--1DONC0#REsCRCD#k0$RLRbNRFsICRRFV.R3RW0H8EVRFRbHMk=0RR8IH0FERVkRF00bkR0IHER
R-0-RE8CRClOHNbDRF0HMRPlFC
83RkRVMHO0F#MROLNDRR5$:hRz)m 1p7e _HkVG;C8R:hRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85E$'H+oEhFR8IFM0RD$'FhI+2R;
RoLCHRM
RHRRV'R$DoCM0<ERR04RE
CMRRRRRCRs0MksRzhqwR;
RCRRD
#CRRRRRCRs#0kDRR:=$R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0F#MROLND;R

RMVkOF0HMOR#NRDL5:$RR)zh p1me_ 7kGVHCR8;hRR:z h)1emp 17_Q th7R2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMOR#NRDL5=$R>,R$
RRRRRRRRRRRRRRRRhRRRR=>0HF_Mo0CChs52
2;RMRC8kRVMHO0F#MROLND;R

RMVkOF0HMOR#NRDL5:$RR)zh p1me_ 7#GVHCR8;hRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58R$H'EohE+RI8FMR0F$F'DI2+h;R
RLHCoMR
RRVRHRD$'C0MoERR<4ER0CRM
RRRRR0sCkRsMhwq1;R
RRDRC#RC
RRRRR#sCkRD0:$=R;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMOR#N;DL
R
RVOkM0MHFRN#OD5LR$RR:z h)1emp #7_VCHG8h;RRz:Rh1) m pe7Q_1t7h 2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRN#OD5LR$>R=R
$,RRRRRRRRRRRRRRRRRRRh=0>RFM_H0CCos25h2R;
R8CMRMVkOF0HMOR#N;DL
R
RVOkM0MHFR_Q#hNCo0CHPRs5NoRR:z h)1emp #7_VCHG8s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRRRHV0XF_jN45sNo5sEo'H2oE2RR='R4'0MEC
RRRRsRRCs0kMsR0k
C;RRRRCCD#
RRRRsRRCs0kMNRVD;#C
RRRR8CMR;HV
CRRMV8Rk0MOHRFMQh#_C0oNH;PC
R
RVOkM0MHFRMVH8H_solE0FR#05oNsRz:Rh1) m pe7V_kH8GC;RR$:aR17p_zmBtQ2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRRV_FsDbFFRV:RFHsRRRHMN'sosCCPs_#CsoNMCFRDFRb
RRRRRRHVN5soH?2R=RR$0MEC
RRRRRRRR0sCkRsMHR;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RsRRCs0kMsRNoH'Eo4E+;RRRRRRRRRRRRRRRR-RR-CRs0MksR0FkRRFVLMFk8'#REEHo
CRRMV8Rk0MOHRFMV8HM_osHEF0l#
0;
VRRk0MOHRFMV8HM_VDC0#lF0NR5s:oRR)zh p1me_ 7kGVHCR8;$RR:1_a7ztpmQ
B2RRRRskC0sQMRhta  H)R#R
RLHCoMR
RRFRVsF_DF:bRRsVFRHHRMsRNoN'sMRoCDbFF
RRRRHRRVsRNo25HRR?=$ER0CRM
RRRRRsRRCs0kM;RH
RRRRCRRMH8RVR;
RCRRMD8RF;Fb
RRRR0sCkRsMN'soD-FI4R;RRRRRRRRRRRRRRRRRRR--skC0sFMRkF0RVFRLk#M8RF'DIR
RCRM8VOkM0MHFRMVH8C_DVF0l#
0;
VRRk0MOHRFMV8HM_osHEF0l#50RNRso:hRz)m 1p7e _H#VG;C8R:$RR71a_mzpt2QB
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RVRRFDs_FRFb:FRVsRRHHNMRsso'CsPC#sC_NCMoRFDFbR
RRRRRHNVRsHo52=R?R0$RE
CMRRRRRRRRskC0sHMR;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RRCRs0MksRoNs'oEHE;+4RRRRRRRRRRRRRRRRR-R-R0sCkRsMFRk0FLVRF8kM#ER'H
oERMRC8kRVMHO0FVMRH_M8sEHo0#lF0
;
RkRVMHO0FVMRH_M8D0CVl0F#Rs5NoRR:z h)1emp #7_VCHG8$;RR1:Raz7_pQmtBR2
RsRRCs0kMhRQa  t)#RH
LRRCMoH
RRRRsVF_FDFbRR:VRFsHMRHRoNs'MsNoDCRF
FbRRRRRVRHRoNs5RH2?$=RRC0EMR
RRRRRRCRs0MksR
H;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRRskC0sNMRsDo'F4I-;RRRRRRRRRRRRRRRRRRR-s-RCs0kMkRF0VRFRkLFMR8#'IDF
CRRMV8Rk0MOHRFMV8HM_VDC0#lF0
;
RkRVMHO0F"MR#"DDR)5qtRR:z h)1emp k7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp z7_ht1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0kF_M5#RN2so;R
RRsRNoP#DRR:=N#soD#PRDBDRmazh;R
RRCRs#0kDRR:=0VF_H8GCRs5NoP#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HM#R"D;D"
R
RVOkM0MHFRs"#D5"RqR)t:hRz)m 1p7e _HkVG;C8RzBmh:aRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDRoNs#RDP:hRz)m 1p7e _1zhQ th7NR5sDo'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58RN'sosoNMC
2;RCRLo
HMRRRRN#soD:PR=FR0_#kMRs5No
2;RRRRN#soD:PR=sRNoP#DRD#sRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"D#s"
;
RkRVMHO0F"MRs"FDR)5qtRR:z h)1emp k7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp z7_ht1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0kF_M5#RN2so;R
RRsRNoP#DRR:=N#soDsPRFBDRmazh;R
RRCRs#0kDRR:=0VF_H8GCRs5NoP#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMsR"F;D"
R
RVOkM0MHFRF"ss5"RqR)t:hRz)m 1p7e _HkVG;C8RzBmh:aRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDRoNs#RDP:hRz)m 1p7e _1zhQ th7NR5sDo'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58RN'sosoNMC
2;RCRLo
HMRRRRN#soD:PR=FR0_#kMRs5No
2;RRRRN#soD:PR=sRNoP#DRssFRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"ssF"
;
RkRVMHO0F"MR#"DNR)5qtRR:z h)1emp k7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp z7_ht1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0kF_M5#RN2so;R
RR-R-RHqs0CEl0RHO#VEH0MRFRRNMkHM#o8MCRRH#NFRDoNHODER#H
V0RRRRN#soD:PR=sRNoP#DRD#DRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"N#D"
;
RkRVMHO0F"MR#"sNR)5qtRR:z h)1emp k7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp z7_ht1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0kF_M5#RN2so;R
RR-R-RHqs0CEl0RHO#VEH0MRFRRNMkHM#o8MCRRH#NFRDoNHODER#H
V0RRRRN#soD:PR=sRNoP#DRD#sRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"N#s"
;
RkRVMHO0F"MR#"DDR)5qtRR:z h)1emp #7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp 17_Q th7NR5sDo'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RN'sosoNMC
2;RCRLo
HMRRRRN#soD:PR=FR0_5#RN2so;R
RRsRNoP#DRR:=N#soD#PRDBDRmazh;R
RRCRs#0kDRR:=0VF_H8GCRs5NoP#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HM#R"D;D"
R
RVOkM0MHFRs"#D5"RqR)t:hRz)m 1p7e _H#VG;C8RzBmh:aRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRPHNsNCLDRoNs#RDP:hRz)m 1p7e _t1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0#F_Rs5No
2;RRRRN#soD:PR=sRNoP#DRD#sRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"D#s"
;
RkRVMHO0F"MRs"FDR)5qtRR:z h)1emp #7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp 17_Q th7NR5sDo'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RN'sosoNMC
2;RCRLo
HMRRRRN#soD:PR=FR0_5#RN2so;R
RRsRNoP#DRR:=N#soDsPRFBDRmazh;R
RRCRs#0kDRR:=0VF_H8GCRs5NoP#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMsR"F;D"
R
RVOkM0MHFRF"ss5"RqR)t:hRz)m 1p7e _H#VG;C8RzBmh:aRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRPHNsNCLDRoNs#RDP:hRz)m 1p7e _t1QhR 75oNs'MDCo-0E4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCRs5NoN'sM2oC;R
RLHCoMR
RRsRNoP#DRR:=0#F_Rs5No
2;RRRRN#soD:PR=sRNoP#DRssFRzBmh
a;RRRRskC#D:0R=FR0_GVHC58RN#soDRP,skC#DE0'H,oER#sCk'D0D2FI;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"ssF"
;
RkRVMHO0F"MR#"DNR)5qtRR:z h)1emp #7_VCHG8B;RmazhRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDNCRsDo#PRR:z h)1emp 17_Q th7NR5sDo'C0MoER-48MFI0jFR2R;
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RN'sosoNMC
2;RCRLo
HMRRRRN#soD:PR=FR0_5#RN2so;R
RRVRHRzBmh>aRR0jRE
CMRRRRR-R-RHqs0CEl0RHO#VEH0CRDVF0RMRRN.R'#ObFlDCClMM0RkClLs#RHRDNRFOoHRH#EVR0
RRRRRoNs#RDP:N=RsDo#PDR#DmRBz;ha
RRRR#CDCR
RRRRRN#soD:PR=sRNoP#DRN#sRm-Bz;ha
RRRR8CMR;HV
RRRR#sCkRD0:0=RFH_VGRC85oNs#,DPR#sCk'D0EEHo,CRs#0kD'IDF2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRD"#N
";
VRRk0MOHRFM"N#s"qR5):tRR)zh p1me_ 7#GVHCR8;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCN#soD:PRR)zh p1me_ 71hQt 57RN'soDoCM04E-RI8FMR0Fj
2;RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85oNs'MsNo;C2
LRRCMoH
RRRRoNs#RDP:0=RFR_#5oNs2R;
RHRRVmRBzRha>RRj0MEC
RRRRNRRsDo#P=R:RoNs#RDP#RsNBhmzaR;
RCRRD
#CRRRRR-R-RHqs0CEl0RHO#VEH0CRDVF0RMRRN.R'#ObFlDCClMM0RkClLs#RHRDNRFOoHRH#EVR0
RRRRRoNs#RDP:N=RsDo#PDR#DBR-mazh;R
RRMRC8VRH;R
RRCRs#0kDRR:=0VF_H8GCRs5NoP#D,CRs#0kD'oEHEs,RCD#k0F'DI
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HM#R"s;N"
R
R-A-RCkON##CRFRlCbbCFDICRNRM00RECFCD8skRVMHO0F3M#
VRRk0MOHRFM1w]Qa _pw5aRqR)t:hRz)m 1p7e _HkVG;C8RzBmh:aRRahqzp)q2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRVRHR)5qtC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwqz;R
RRMRC8VRH;R
RRCRs0MksRtq)RN#DRzBmh
a;RMRC8kRVMHO0F1MR]aQw_wp a
;
RkRVMHO0F1MR]aQw_t)Q]5aRqR)t:hRz)m 1p7e _HkVG;C8RzBmh:aRRahqzp)q2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRVRHR)5qtC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwqz;R
RRMRC8VRH;R
RRCRs0MksRtq)RN#sRzBmh
a;RMRC8kRVMHO0F1MR]aQw_t)Q]
a;
VRRk0MOHRFM1w]Qa _pw5aRqR)t:hRz)m 1p7e _H#VG;C8RzBmh:aRRahqzp)q2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRVRHR)5qtC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRCRs0MksRtq)RN#DRzBmh
a;RMRC8kRVMHO0F1MR]aQw_wp a
;
RkRVMHO0F1MR]aQw_t)Q]5aRqR)t:hRz)m 1p7e _H#VG;C8RzBmh:aRRahqzp)q2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRVRHR)5qtC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRCRs0MksRtq)RN#sRzBmh
a;RMRC8kRVMHO0F1MR]aQw_t)Q]
a;
-RR-------------------------------------------------------------------------
--R-R-RoDFHDONRMVkOF0HMR#
R----------------------------------------------------------------------------R
RVOkM0MHFRF"M05"RpRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RR R)1azpRR:=MRF00#F_k5DPp
2;RRRRskC0s0MRFV_kH8GC51) z,paREp'H,oERDp'F;I2
CRRMV8Rk0MOHRFM"0MF"
;
RkRVMHO0F"MRN"M8R,5pR:)RR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52MRN8FR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"N""M"8":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0kF_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM""FsR,5pR:)RR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52sRFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"s"F"R":)oNMCsRCsRFspq')hRt /)=R'h)qt
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRR)z 1p:aR=FR50sEC#>R=R''X2R;
RCRRMH8RVR;
RsRRCs0kMFR0_HkVG5C8)z 1pRa,pH'EoRE,pF'DI
2;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRN"MMR8"5Rp,)RR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRMMN8FR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"M""N"M8"):RNCMoRsCsFpsR'h)qt/ R='R))tqh R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRR)RR p1za=R:R05FE#CsRR=>'2X';R
RRMRC8VRH;R
RRCRs0MksR_0FkGVHC)85 p1zap,R'oEHEp,R'IDF2R;
R8CMRMVkOF0HMMR"N"M8;R

RMVkOF0HMMR"FRs"5Rp,)RR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRsMFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"F"Ms:""RM)NoCCRsssFR)p'q htRR/=)q')h"t 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR1) zRpa:5=RFC0Es=#R>XR''
2;RRRRCRM8H
V;RRRRskC0s0MRFV_kH8GC51) z,paREp'H,oERDp'F;I2
CRRMV8Rk0MOHRFM"sMF"
;
RkRVMHO0F"MRG"FsR,5pR:)RR)zh p1me_ 7kGVHCR82skC0szMRh1) m pe7V_kH8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52FRGsFR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"G""F"s":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0kF_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"Rp),RRz:Rh1) m pe7V_kH8GC2CRs0MksR)zh p1me_ 7kGVHCH8R#R
RRNRPsLHND)CR p1zaRR:1_a7ztpmQeB_ mBa)'5pDoCM04E-RI8FMR0FjR2;RR--VOFsCFR8IFM0
LRRCMoH
RRRRRHV5Ep'HRoE='R)EEHoR8NMRDp'F=IRRD)'FRI20MEC
RRRR)RR p1za=R:R_0F#PkD5Rp2GsMFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"M"GF"s":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0kF_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRM"GF;s"
R
RVOkM0MHFRF"M05"RpRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RR R)1azpRR:=MRF00#F_k5DPp
2;RRRRskC0s0MRFV_#H8GC51) z,paREp'H,oERDp'F;I2
CRRMV8Rk0MOHRFM"0MF"
;
RkRVMHO0F"MRN"M8R,5pR:)RR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52MRN8FR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"N""M"8":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0#F_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM""FsR,5pR:)RR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52sRFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"s"F"R":)oNMCsRCsRFspq')hRt /)=R'h)qt
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRR)z 1p:aR=FR50sEC#>R=R''X2R;
RCRRMH8RVR;
RsRRCs0kMFR0_H#VG5C8)z 1pRa,pH'EoRE,pF'DI
2;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRN"MMR8"5Rp,)RR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRMMN8FR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"M""N"M8"):RNCMoRsCsFpsR'h)qt/ R='R))tqh R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRR)RR p1za=R:R05FE#CsRR=>'2X';R
RRMRC8VRH;R
RRCRs0MksR_0F#GVHC)85 p1zap,R'oEHEp,R'IDF2R;
R8CMRMVkOF0HMMR"N"M8;R

RMVkOF0HMMR"FRs"5Rp,)RR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VGRC8HR#
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmp)5'MDCo-0E4FR8IFM0R;j2R-R-RsVFO8CRF0IMFR
RLHCoMR
RRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRsMFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"F"Ms:""RM)NoCCRsssFR)p'q htRR/=)q')h"t 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR1) zRpa:5=RFC0Es=#R>XR''
2;RRRRCRM8H
V;RRRRskC0s0MRFV_#H8GC51) z,paREp'H,oERDp'F;I2
CRRMV8Rk0MOHRFM"sMF"
;
RkRVMHO0F"MRG"FsR,5pR:)RR)zh p1me_ 7#GVHCR82skC0szMRh1) m pe7V_#H8GCR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RHRRVpR5'oEHERR=)H'EoNERMp8R'IDFR)=R'IDF2ER0CRM
RRRRR1) zRpa:0=RFk_#DpP52FRGsFR0_D#kP25);R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"G""F"s":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0#F_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"Rp),RRz:Rh1) m pe7V_#H8GC2CRs0MksR)zh p1me_ 7#GVHCH8R#R
RRNRPsLHND)CR p1zaRR:1_a7ztpmQeB_ mBa)'5pDoCM04E-RI8FMR0FjR2;RR--VOFsCFR8IFM0
LRRCMoH
RRRRRHV5Ep'HRoE='R)EEHoR8NMRDp'F=IRRD)'FRI20MEC
RRRR)RR p1za=R:R_0F#PkD5Rp2GsMFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"M"GF"s":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0#F_VCHG8 5)1azp,'RpEEHo,'RpD2FI;R
RCRM8VOkM0MHFRM"GF;s"
R
R-e-RCFO0sMRN80R#8D_kFOoHRMVkOF0HMR#,#CNlRRN#VOkM0MHF#MRHRlMkCOsH_8#0
VRRk0MOHRFM"8NM"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85s)'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RNpRM)8R5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7V_kH8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52MRN8;R)
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM""FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58R)N'sM2oC;R
RLHCoMR
RRFRVsRRHHsMRCD#k0N'sMRoCDbFF
RRRRsRRCD#k025HRR:=psRFRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRs"F"pR5Rz:Rh1) m pe7V_kH8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52sRFR
);RRRRCRM8DbFF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM""Fs;R

RMVkOF0HMMR"N"M8RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58R)N'sM2oC;R
RLHCoMR
RRFRVsRRHHsMRCD#k0N'sMRoCDbFF
RRRRsRRCD#k025HRR:=pNRMM)8R5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRN"MM;8"
R
RVOkM0MHFRN"MMR8"5:pRR)zh p1me_ 7kGVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp k7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2M8NMR
);RRRRCRM8DbFF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"MMN8
";
VRRk0MOHRFM"sMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85s)'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RMpRF)sR5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Ms
";
VRRk0MOHRFM"sMF"pR5Rz:Rh1) m pe7V_kH8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52FRMs;R)
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Ms
";
VRRk0MOHRFM"sGF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85s)'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RGpRF)sR5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7V_kH8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52FRGs;R)
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"RpRR:1_a7ztpmQRB;)RR:z h)1emp k7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCR'5)soNMC
2;RCRLo
HMRRRRVRFsHMRHR#sCk'D0soNMCFRDFRb
RRRRR#sCk5D0H:2R=RRpGsMFRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRGsMF"
;
RkRVMHO0F"MRGsMF"pR5Rz:Rh1) m pe7V_kH8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52MRGF)sR;R
RRMRC8FRDF
b;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMGR"M"Fs;R

RMVkOF0HMNR"MR8"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8)R5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=RR8NMRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRN"M8;R

RMVkOF0HMNR"MR8"5:pRR)zh p1me_ 7#GVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2NRM8)R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRN"M8;R

RMVkOF0HMFR"s5"RpRR:1_a7ztpmQRB;)RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCR'5)soNMC
2;RCRLo
HMRRRRVRFsHMRHR#sCk'D0soNMCFRDFRb
RRRRR#sCk5D0H:2R=RRpF)sR5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRs"F"
;
RkRVMHO0F"MRFRs"5:pRR)zh p1me_ 7#GVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2F)sR;R
RRMRC8FRDF
b;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFR"s
";
VRRk0MOHRFM"MMN85"RpRR:1_a7ztpmQRB;)RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCR'5)soNMC
2;RCRLo
HMRRRRVRFsHMRHR#sCk'D0soNMCFRDFRb
RRRRR#sCk5D0H:2R=RRpM8NMRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRM8NM"
;
RkRVMHO0F"MRM8NM"pR5Rz:Rh1) m pe7V_#H8GC;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85sp'NCMo2R;
RoLCHRM
RVRRFHsRRRHMskC#Ds0'NCMoRFDFbR
RRRRRskC#DH052=R:RHp52NRMM)8R;R
RRMRC8FRDF
b;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMMR"N"M8;R

RMVkOF0HMMR"FRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8)R5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=RRsMFRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRM"Fs;R

RMVkOF0HMMR"FRs"5:pRR)zh p1me_ 7#GVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2MRFs)R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRM"Fs;R

RMVkOF0HMGR"FRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8)R5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=RRsGFRH)52R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRG"Fs;R

RMVkOF0HMGR"FRs"5:pRR)zh p1me_ 7#GVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2GRFs)R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRG"Fs;R

RMVkOF0HMGR"M"FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _H#VG2C8
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58R)N'sM2oC;R
RLHCoMR
RRFRVsRRHHsMRCD#k0N'sMRoCDbFF
RRRRsRRCD#k025HRR:=pMRGF)sR5;H2
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRM"GF;s"
R
RVOkM0MHFRM"GFRs"5:pRR)zh p1me_ 7#GVHCR8;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8pR5'MsNo;C2
LRRCMoH
RRRRsVFRHHRMCRs#0kD'MsNoDCRF
FbRRRRRCRs#0kD5RH2:p=R5RH2GsMFR
);RRRRCRM8DbFF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"FGMs
";
-RR-CR)80kOHRFMFsbCNs0F#R
RVOkM0MHFRM"N85"RDRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sNMRM08RFk_#DDP52R;
R8CMRMVkOF0HMNR"M;8"
R
RVOkM0MHFRN"MMR8"5:DRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMM8NMR_0F#PkD5;D2
CRRMV8Rk0MOHRFM"MMN8
";
VRRk0MOHRFM""FsRR5D:hRz)m 1p7e _HkVG2C8R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRRFs0#F_k5DPD
2;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRF"Ms5"RDRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sMMRF0sRFk_#DDP52R;
R8CMRMVkOF0HMMR"F;s"
R
RVOkM0MHFRF"Gs5"RDRR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sGMRF0sRFk_#DDP52R;
R8CMRMVkOF0HMGR"F;s"
R
RVOkM0MHFRM"GFRs"5:DRR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMGsMFR_0F#PkD5;D2
CRRMV8Rk0MOHRFM"FGMs
";
VRRk0MOHRFM"8NM"DR5Rz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMMRN8FR0_D#kP25D;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM"MMN85"RDRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sMMRNRM80#F_k5DPD
2;RMRC8kRVMHO0F"MRM8NM"
;
RkRVMHO0F"MRFRs"5:DRR)zh p1me_ 7#GVHCR82skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMF0sRFk_#DDP52R;
R8CMRMVkOF0HMFR"s
";
VRRk0MOHRFM"sMF"DR5Rz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMFRMsFR0_D#kP25D;R
RCRM8VOkM0MHFRF"Ms
";
VRRk0MOHRFM"sGF"DR5Rz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMFRGsFR0_D#kP25D;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"RDRR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sGMRMRFs0#F_k5DPD
2;RMRC8kRVMHO0F"MRGsMF"R;
RR-- RM8skC8OF0HMbRFC0sNF
s#
VRRk0MOHRFM""?=R,5pR:)RR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo;E2
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=l#HM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCDP#D,#RsDRPRRRRRRz:Rh1) m pe7h_z1hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RCRLoRHMRR--?R=
RHRRV5R5pC'DMEo0R4<R2sRFR'5)DoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"="?"R":MDkDR08CCCO08s,RCs0kMoHMR
X"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s'MRX
';RRRRCCD#
RRRRDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRCss#CHxRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDRR#RDPR:RR=FR0_#kMRs5DCx#HC
2;RRRRR#RsDRPRR=R:R_0FkRM#5Css#CHx2R;
RRRRR0sCkRsMDP#DRR?=sP#D;R
RRMRC8VRH;R
RCRM8VOkM0MHFR="?"
;
RkRVMHO0F"MR?"/=R,5pR:)RR)zh p1me_ 7kGVHCR82skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo;E2
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=l#HM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCDP#D,#RsDRPRRRRRRz:Rh1) m pe7h_z1hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RCRLoRHMRR--?
/=RRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"?""/"=":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRR:=0kF_M5#RD#sCH2xC;R
RRRRRsP#DRRRR:0=RFM_k#sR5sHC#x;C2
RRRRsRRCs0kM#RDD?PR/s=R#;DP
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?/"
;
RkRVMHO0F"MR?R>"5Rp,)RR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _1zhQ th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRMR-?-R>R
RRVRHRD55'MDCoR0E<2R4RRFs5Ds'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""?>"M:RkRDD8CC0O80C,CRs0MksHRMoXR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRR#RDDRPRR=R:R_0FkRM#5CDs#CHx2R;
RRRRRDs#PRRRRR:=0kF_M5#Rs#sCH2xC;R
RRRRRskC0sDMR#RDP?s>R#;DP
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?>;R

RMVkOF0HM?R">R="5Rp,)RR:z h)1emp k7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _1zhQ th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRMR-?-R>R=
RHRRV5R5DC'DMEo0R4<R2sRFR'5sDoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R">"?=:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRDP#DRRRR:0=RFM_k#DR5sHC#x;C2
RRRRsRR#RDPR:RR=FR0_#kMRs5sCx#HC
2;RRRRRCRs0MksRDD#P>R?=#RsD
P;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<5"Rp),RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLC#RDDRP,sP#DRRRRR:RRR)zh p1me_ 7zQh1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoM-RR-<R?
RRRRRHV5'5DDoCM0<ERRR42F5sRsC'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""?"<":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRR:=0kF_M5#RD#sCH2xC;R
RRRRRsP#DRRRR:0=RFM_k#sR5sHC#x;C2
RRRRsRRCs0kM#RDD?PR<#RsD
P;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;<"
R
RVOkM0MHFR<"?=5"Rp),RRz:Rh1) m pe7V_kH8GC2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLC#RDDRP,sP#DRRRRR:RRR)zh p1me_ 7zQh1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoM-RR-<R?=R
RRVRHRD55'MDCoR0E<2R4RRFs5Ds'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""=?<"R":MDkDR08CCCO08s,RCs0kMoHMR
X"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s'MRX
';RRRRCCD#
RRRRDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRCss#CHxRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDRR#RDPR:RR=FR0_#kMRs5DCx#HC
2;RRRRR#RsDRPRR=R:R_0FkRM#5Css#CHx2R;
RRRRR0sCkRsMDP#DR=?<RDs#PR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
RVOkM0MHFR="?"pR5,RR):hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQHBR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRMR-?-R=R
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""?="M:RkRDD8CC0O80C,CRs0MksHRMoXR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRR#RDDRPRR=R:R_0F#DR5sHC#x;C2
RRRRsRR#RDPR:RR=FR0_5#Rs#sCH2xC;R
RRRRRskC0sDMR#RDP?s=R#;DP
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?=;R

RMVkOF0HM?R"/R="5Rp,)RR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _t1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoHR-R-R=?/
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""?"/="M:RkRDD8CC0O80C,CRs0MksHRMoXR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRR#RDDRPRR=R:R_0F#DR5sHC#x;C2
RRRRsRR#RDPR:RR=FR0_5#Rs#sCH2xC;R
RRRRRskC0sDMR#RDP?R/=sP#D;R
RRMRC8VRH;R
RCRM8VOkM0MHFR/"?=
";
VRRk0MOHRFM""?>R,5pR:)RR)zh p1me_ 7#GVHCR82skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo;E2
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=l#HM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp #7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCDP#D,#RsDRPRRRRRRz:Rh1) m pe7Q_1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoM-RR->R?
RRRRRHV5'5DDoCM0<ERRR42F5sRsC'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""?">":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRR:=0#F_Rs5DCx#HC
2;RRRRR#RsDRPRR=R:R_0F#sR5sHC#x;C2
RRRRsRRCs0kM#RDD?PR>#RsD
P;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;>"
R
RVOkM0MHFR>"?=5"Rp),RRz:Rh1) m pe7V_#H8GC2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLC#RDDRP,sP#DRRRRR:RRR)zh p1me_ 71hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RCRLoRHMRR--?
>=RRRRH5VR5DD'C0MoERR<4F2RssR5'MDCoR0E<2R42ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"?"">"=":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RRRRRDD#PRRRRR:=0#F_Rs5DCx#HC
2;RRRRR#RsDRPRR=R:R_0F#sR5sHC#x;C2
RRRRsRRCs0kM#RDD?PR>s=R#;DP
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?>"
;
RkRVMHO0F"MR?R<"5Rp,)RR:z h)1emp #7_VCHG8s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _t1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoHR-R-R
?<RRRRH5VR5DD'C0MoERR<4F2RssR5'MDCoR0E<2R42ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"?""<:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRDP#DRRRR:0=RFR_#5CDs#CHx2R;
RRRRRDs#PRRRRR:=0#F_Rs5sCx#HC
2;RRRRRCRs0MksRDD#P<R?RDs#PR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
VRRk0MOHRFM"=?<"pR5,RR):hRz)m 1p7e _H#VG2C8R0sCkRsM1_a7ztpmQHBR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRMR-?-R<R=
RHRRV5R5DC'DMEo0R4<R2sRFR'5sDoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"<"?=:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RRRRRDP#DRRRR:0=RFR_#5CDs#CHx2R;
RRRRRDs#PRRRRR:=0#F_Rs5sCx#HC
2;RRRRRCRs0MksRDD#P<R?=#RsD
P;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?"<=;R

RR--vON0EkRVMHO0FRM,#HHlDRNs0"FR#_08lON0EV"RsRFlMCkls_HO#
08RkRVMHO0F#MR0l8_NE0OR,5pR:)RR)zh p1me_ 7kGVHCR82skC0sAMRm mpqHhR#R
RLHCoMR
RRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRRskC0s#MR0l8_NE0O5_0F#PkD5,p2R_0F#PkD52)2;R
RRDRC#RC
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"71a_avqBR]:pq')hRt /)=R'h)qtR ,skC0sMMHoqRwp"1 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMV#NDCR;
RCRRMH8RVR;
R8CMRMVkOF0HM0R#8N_l0;OE
R
RVOkM0MHFR8#0_0lNO5ERp),RRz:Rh1) m pe7V_#H8GC2CRs0MksRmAmph qR
H#RCRLo
HMRRRRH5VRpH'Eo=ERRE)'HRoENRM8pF'DIRR=)F'DI02RE
CMRRRRRCRs0MksR8#0_0lNO0E5Fk_#DpP520,RFk_#D)P52
2;RRRRCCD#
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&1R"av7_q]aB:'Rp)tqh =R/R))'q ht,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR8CMR;HV
CRRMV8Rk0MOHRFM#_08lON0E
;
R-R-RlOFbCNsRMVkOF0HMR#
RMVkOF0HM=R""
R5RRRRDs,RRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm 
qhR#RH
RRRRMOF#M0N0CRDVH0_MG8CRRRRR:RRRaQh )t RR:=lHNGl5klDH'EoRE,sH'Eo;E2
RRRRMOF#M0N0HRso_E0HCM8GRRRR:RRRaQh )t RR:=l#HM5DD'FRI,sF'DI
2;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCDP#D,#RsDRPRRRRRRz:Rh1) m pe7h_z1hQt 57RD#sCH'xCDoCM04E-RI8FMR0Fj
2;RCRLo
HMRRRRH5VRDC'DMEo0R4<RRRFssC'DMEo0R4<R2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"="""R":MDkDRoNskMlC0CR800COCR8,skC0sMMHoqRwp"1 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMV#NDCR;
RCRRDV#HR#5Q_DX52sRFR_Q#X25s2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"="""R":lNC0PkNDCCR800COCR8,skC0sMMHoqRwp"1 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMV#NDCR;
RCRRMH8RVR;
RDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RDRR#RDPR:RR=FR0_#kMRs5DCx#HC
2;RRRRsP#DRRRR:0=RFM_k#sR5sHC#x;C2
RRRR0sCkRsMDP#DRs=R#;DP
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR""=RR5
RDRR,RRs:hRz)m 1p7e _H#VG2C8RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqRh
R
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _t1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""=:""RDMkDsRNoCklM80RCO0C0,C8R0sCkHsMMwoRq p1"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRDVN#
C;RRRRCHD#VQR5#5_XDF2Rs#RQ_sX5202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""=:""R0lCNDPNk8CRCO0C0,C8R0sCkHsMMwoRq p1"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRDVN#
C;RRRRCRM8H
V;RRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRDP#DRRRR:0=RFR_#5CDs#CHx2R;
RsRR#RDPR:RR=FR0_5#Rs#sCH2xC;R
RRCRs0MksRDD#PRR=sP#D;R
RCRM8VOkM0MHFR""=;R

RMVkOF0HM/R"=5"R
RRRRRD,sRR:z h)1emp k7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp z7_ht1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""/"=":kRMDNDRslokCRM08CC0O80C,CRs0MksHRMoa )z"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRk0sCR;
RCRRDV#HR#5Q_DX52sRFR_Q#X25s2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"/""=:""R0lCNDPNk8CRCO0C0,C8R0sCkHsMMaoR)"z 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM0Csk;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RR#RDDRPRR=R:R_0FkRM#5CDs#CHx2R;
RsRR#RDPR:RR=FR0_#kMRs5sCx#HC
2;RRRRskC0sDMR#RDP/s=R#;DP
CRRMV8Rk0MOHRFM""/=;R

RMVkOF0HM/R"=5"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"="/"R":MDkDRoNskMlC0CR800COCR8,skC0sMMHo)Raz
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s0MRs;kC
RRRR#CDH5VRQX#_5RD2FQsR#5_XsR220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""/="l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRza) R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMsR0k
C;RRRRCRM8H
V;RRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRDP#DRRRR:0=RFR_#5CDs#CHx2R;
RsRR#RDPR:RR=FR0_5#Rs#sCH2xC;R
RRCRs0MksRDD#P=R/RDs#PR;
R8CMRMVkOF0HM/R"=
";
VRRk0MOHRFM"R>"5R
RR,RDR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp hR
RHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLC#RDDRP,sP#DRRRRR:RRR)zh p1me_ 7zQh1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRR420MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""">":kRMDNDRslokCRM08CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR#CDH5VRQX#_5RD2FQsR#5_XsR220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""">":CRl0NNPDRkC8CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR8CMR;HV
RRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRCss#CHxRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDD#PRRRRR:=0kF_M5#RD#sCH2xC;R
RR#RsDRPRR=R:R_0FkRM#5Css#CHx2R;
RsRRCs0kM#RDD>PRRDs#PR;
R8CMRMVkOF0HM>R""
;
RkRVMHO0F"MR>5"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R""">"M:RkRDDNksol0CMR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRDRC#RHV5_Q#X25DRRFsQX#_52s2RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R""">"l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RR#RDDRPRR=R:R_0F#DR5sHC#x;C2
RRRRDs#PRRRRR:=0#F_Rs5sCx#HC
2;RRRRskC0sDMR#RDP>#RsD
P;RMRC8kRVMHO0F"MR>
";
VRRk0MOHRFM"R<"5R
RR,RDR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp hR
RHR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRsPNHDNLC#RDDRP,sP#DRRRRR:RRR)zh p1me_ 7zQh1t7h Rs5DCx#HCC'DMEo0-84RF0IMF2Rj;R
RLHCoMR
RRVRHR'5DDoCM0<ERRF4Rs'RsDoCM0<ERRR420MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""<":kRMDNDRslokCRM08CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR#CDH5VRQX#_5RD2FQsR#5_XsR220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""<":CRl0NNPDRkC8CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR8CMR;HV
RRRRCDs#CHxRR:=sHC#x5CRDD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRCss#CHxRR:=sHC#x5CRsD,RC_V0HCM8Gs,RH0oE_8HMC;G2
RRRRDD#PRRRRR:=0kF_M5#RD#sCH2xC;R
RR#RsDRPRR=R:R_0FkRM#5Css#CHx2R;
RsRRCs0kM#RDD<PRRDs#PR;
R8CMRMVkOF0HM<R""
;
RkRVMHO0F"MR<5"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"""<"M:RkRDDNksol0CMR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRDRC#RHV5_Q#X25DRRFsQX#_52s2RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"""<"l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RR#RDDRPRR=R:R_0F#DR5sHC#x;C2
RRRRDs#PRRRRR:=0#F_Rs5sCx#HC
2;RRRRskC0sDMR#RDP<#RsD
P;RMRC8kRVMHO0F"MR<
";
VRRk0MOHRFM"">=RR5
RDRR,RRs:hRz)m 1p7e _HkVG2C8RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqRh
R
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _1zhQ th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"=">"R":MDkDRoNskMlC0CR800COCR8,skC0sMMHoqRwp"1 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMV#NDCR;
RCRRDV#HR#5Q_DX52sRFR_Q#X25s2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&">""=:""R0lCNDPNk8CRCO0C0,C8R0sCkHsMMwoRq p1"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRDVN#
C;RRRRCRM8H
V;RRRRD#sCHRxC:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxC:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRDP#DRRRR:0=RFM_k#DR5sHC#x;C2
RRRRDs#PRRRRR:=0kF_M5#Rs#sCH2xC;R
RRCRs0MksRDD#P=R>RDs#PR;
R8CMRMVkOF0HM>R"=
";
VRRk0MOHRFM"">=RR5
RDRR,RRs:hRz)m 1p7e _H#VG2C8RRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqRh
R
H#RRRRO#FM00NMRVDC0M_H8RCGRRRRRRR:Q hatR ):l=RNlGHkDl5'oEHEs,R'oEHE
2;RRRRO#FM00NMRosHEH0_MG8CRRRRRRR:Q hatR ):l=RH5M#DF'DIs,R'IDF2R;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDDCR#,DPRDs#PRRRRRRR:hRz)m 1p7e _t1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR""">"=":kRMDNDRslokCRM08CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR#CDH5VRQX#_5RD2FQsR#5_XsR220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""">="l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RRsRDCx#HC=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HC=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RR#RDDRPRR=R:R_0F#DR5sHC#x;C2
RRRRDs#PRRRRR:=0#F_Rs5sCx#HC
2;RRRRskC0sDMR#RDP>s=R#;DP
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"R
RRRRRD,sRR:z h)1emp k7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp z7_ht1QhR 75CDs#CHx'MDCo-0E4FR8IFM0R;j2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRR"""<"=":kRMDNDRslokCRM08CC0O80C,CRs0MksHRMow1qp R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMNRVD;#C
RRRR#CDH5VRQX#_5RD2FQsR#5_XsR220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""<="l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRpwq1
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RRsRDCx#HCRRRR=R:R#sCHRxC5RD,D0CV_8HMCRG,sEHo0M_H82CG;R
RRsRsCx#HCRRRR=R:R#sCHRxC5Rs,D0CV_8HMCRG,sEHo0M_H82CG;R
RR#RDDRPRRRRRR=R:R_0FkRM#5CDs#CHx2R;
RsRR#RDPRRRRR:RR=FR0_#kMRs5sCx#HC
2;RRRRskC0sDMR#RDP<s=R#;DP
CRRMV8Rk0MOHRFM""<=;R

RMVkOF0HM<R"=5"R
RRRRRD,sRR:z h)1emp #7_VCHG8R2RRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MD0RC_V0HCM8GRRRRRRR:hRQa  t)=R:RGlNHllk5ED'H,oEREs'H2oE;R
RRFROMN#0Ms0RH0oE_8HMCRGRRRRR:hRQa  t)=R:RMlH#'5DD,FIRDs'F;I2
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRDD#Ps,R#RDPRRRRRRR:z h)1emp 17_Q th7DR5sHC#xDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVDR5'MDCoR0E<RR4FssR'MDCoR0E<2R4RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"="<"R":MDkDRoNskMlC0CR800COCR8,skC0sMMHoqRwp"1 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMV#NDCR;
RCRRDV#HR#5Q_DX52sRFR_Q#X25s2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"<""=:""R0lCNDPNk8CRCO0C0,C8R0sCkHsMMwoRq p1"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRDVN#
C;RRRRCRM8H
V;RRRRD#sCHRxCRRRR:s=RCx#HCDR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRs#sCHRxCRRRR:s=RCx#HCsR5,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRDP#DRRRRRRRR:0=RFR_#5CDs#CHx2R;
RsRR#RDPRRRRR:RR=FR0_5#Rs#sCH2xC;R
RRCRs0MksRDD#P=R<RDs#PR;
R8CMRMVkOF0HM<R"=
";
-RR-PRFCFsDNR8#F0VRE8CRCkVNDl0RNlGHkNlRMl8RHlMHkVlRk0MOH#FM
VRRk0MOHRFMlHNGlRkl5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVGRC8HR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMFR0_GVHCl85NlGHk0l5FM_k#s5DCx#HCR2,0kF_Ms#5sHC#x2C2,R
RRRRRRRRRRRRRRRRRRCRDVH0_MG8C,HRso_E0HCM8G
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHNGlRkl5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VGRC8HR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMFR0_GVHCl85NlGHk0l5F5_#D#sCH2xC,FR0_s#5sHC#x2C2,R
RRRRRRRRRRRRRRRRRRCRDVH0_MG8C,HRso_E0HCM8G
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5RD,sRR:z h)1emp k7_VCHG8s2RCs0kMhRz)m 1p7e _HkVGRC8HR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMFR0_GVHCl85HlMHk0l5FM_k#s5DCx#HCR2,0kF_Ms#5sHC#x2C2,R
RRRRRRRRRRRRRRRRRRCRDVH0_MG8C,HRso_E0HCM8G
2;RMRC8kRVMHO0FlMRHlMHk
l;
VRRk0MOHRFMlHHMlRkl5RD,sRR:z h)1emp #7_VCHG8s2RCs0kMhRz)m 1p7e _H#VGRC8HR#
RORRF0M#NRM0D0CV_8HMCRGRRRRRRQ:Rhta  :)R=NRlGkHll'5DEEHo,'RsEEHo2R;
RORRF0M#NRM0sEHo0M_H8RCGRRRRRQ:Rhta  :)R=HRlMD#5'IDF,'RsD2FI;R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
LRRCMoH
RRRRRHV5DD'C0MoERR<4sRFRDs'C0MoERR<402RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RDRRsHC#x:CR=CRs#CHxR,5DRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRsHC#x:CR=CRs#CHxR,5sRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMFR0_GVHCl85HlMHk0l5F5_#D#sCH2xC,FR0_s#5sHC#x2C2,R
RRRRRRRRRRRRRRRRRRCRDVH0_MG8C,HRso_E0HCM8G
2;RMRC8kRVMHO0FlMRHlMHk
l;
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:qRhaqz)pR;R-H-RMo0CCRs
RORRF0M#NRM0D0CV_8HMCRGRR:RRRaQh )t ;-RR-CRDVH0RMG8CRH5EoHERMG8C2R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hatR )RRRRRRRRRRRRRRRRR=R:RRj;RR--sEHo0MRH8
CGRRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRMOF#M0N0IRVRRRRRRR:Q hatR ):l=RHRM#5osHEH0_MG8C,HRso_E0HCM8GR2;RR--OON0EHRD0NCsDR#
RPRRNNsHLRDCskC#DR0R:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0VFRI
2;RRRRPHNsNCLDRC#s#0kDRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0Fj:2R=R
RRRRR5EF0CRs#='>Rj;'2R-R-R0HMCsoCRsbF0MHF
RRRRsPNHDNLCsRNoRGRRRR:hzqa);qpRRRRRRRRRR--HCM0sDMNRsPC#MHFRRFVN
soRCRLo
HMRRRRH5VRskC#DD0'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RHRRVsRNo=R/R0jRE
CMRRRRRsRNo:GR=sRNoR;
RRRRRsVFRHQRMRRj0#FRskC#DD0'CRV0DbFF
RRRRRRRRRHV5oNsGFRl82R.Rj=RRC0EMR
RRRRRRRRR##sCk5D0Q:2R=jR''R;
RRRRRCRRD
#CRRRRRRRRRsR#CD#k025QRR:=';4'
RRRRRRRR8CMR;HV
RRRRRRRRoNsG=R:RoNsG;/.
RRRRCRRMD8RF;Fb
RRRRHRRVsRNo/GR=RRj0MEC
RRRRRRRR#N#CRs0hWm_qQ)hhRt
RRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRRRRR&"_amzXwQ h75q)azq:p2ROPC0RFs0MskOCN08R"
RRRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRRHRRVPRFCDsVF#I_0C$DRV=RH8GC_0#Nk0sNCER0CRM
RRRRRRRRR0sCkRsM#kN0sCN0RC5DVH0_MG8C,HRso_E0HCM8G
2;RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRRRRskC#D:0R=CRs#CHxRs5NoRRRRRRRRRRRRR=>##sCk,D0
RRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=D>RC_V0HCM8GR,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=RosHEH0_MG8C,R
RRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRCCD#
RRRRsRRCD#k0=R:R05FE#CsRR=>'2j';R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0kF_VCHG8
;
RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRaQh )t ;-RR-MRH0CCosR
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )R-R-RVDC0MRH8RCG5oEHEMRH82CG
RRRRMOF#M0N0HRso_E0HCM8GRRRRQ:Rhta  R)RRRRRRRRRRRRRRRRRRR:=jR;R-s-RH0oER8HMCRG
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRO#FM00NMRRVIRRRRRQ:Rhta  :)R=HRlM5#RsEHo0M_H8,CGRosHEH0_MG8C2R;R-O-RNE0OR0DHCDsN#R
RRNRPsLHNDsCRCD#k0:RRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFIRV2R;
RPRRNNsHLRDC##sCkRD0:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0jFR2=R:
RRRR5RRFC0Es=#R>jR''R2;RR--HCM0oRCsb0FsH
FMRRRRPHNsNCLDRoNsGRRRRQ:Rhta  R);RRRRRRRR-H-RMs0CMRNDP#CsHRFMFNVRsRo
RPRRNNsHLRDC#MHoRRRR:aR17p_zmBtQ;RRRR-RR-HR#oFMRVMRHb
k0RCRLo
HMRRRRH5VRskC#DD0'C0MoERR<402RERCMRRRRRRRR-M-RkRDDsoNMCR
RRRRRskC0shMRq;1w
RRRR8CMR;HV
RRRRRHVNRso/j=RRC0EMR
RRRRRH5VRNRso<2RjRC0EMR
RRRRRRHR#o:MR=4R''R;
RRRRRNRRsRoG:-=R5oNsR4+R2R;
RRRRR#CDCR
RRRRRRHR#o:MR=jR''R;
RRRRRNRRsRoG:N=Rs
o;RRRRRMRC8VRH;R
RRRRRVRFsQMRHR0jRFsR#CD#k0C'DVD0RF
FbRRRRRRRRH5VRNGsoR8lFRR.2=RRj0MEC
RRRRRRRR#RRskC#DQ052=R:Ro#HMR;
RRRRRCRRD
#CRRRRRRRRRsR#CD#k025QRR:=MRF0#MHo;R
RRRRRRMRC8VRH;R
RRRRRRsRNo:GR=sRNo.G/;R
RRRRRCRM8DbFF;R
RRRRRHNVRsRoG/j=RRRFsD0CV_8HMC<GRRFjRsHR#o/MR=sR#CD#k0s5#CD#k0C'DVR020MEC
RRRRRRRR#N#CRs0hWm_qQ)hhRt
RRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRRRRR&"_am1XwQ Q75hta  :)2ROPC0RFs0MskOCN08R"
RRRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRRHRRVPRFCDsVF#I_0C$DRV=RH8GC_0#Nk0sNCER0CRMRRRRRRRRRRRRRR-R-R0#Nk0sNCR
RRRRRRRRRHNVRs<oRR0jRE
CMRRRRRRRRRRRRskC#D:0R=FRM0NR#0Nks05CRskC#DE0'H,oER#sCk'D0D2FI;-RR-MRk8VCsD
FIRRRRRRRRRDRC#RC
RRRRRRRRRsRRCD#k0=R:R0#Nk0sNCsR5CD#k0H'EoRE,skC#DD0'F;I2RRRRR-R-RCFPsFVDIR
RRRRRRRRRCRM8H
V;RRRRRRRRRCRs0MksR#sCk;D0
RRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RRRRR#sCkRD0:s=RCx#HCNR5sRoRRRRRRRRRR>R=RC#s#0kD,R
RRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>D0CV_8HMC
G,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>HRso_E0HCM8GR,
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRR#CDCR
RRRRRskC#D:0R=FR50sEC#>R=R''j2R;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0F#GVHC
8;
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)qRp;RRRR-s-RC
NDRRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-D-RCRV0HCM8GER5HRoEHCM8GR2
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;-RR-HRsoRE0HCM8GR
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02-RR-RRyFoVRk8NsR0LH#R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMRRVIRRRRRRRRRRRRRQ:Rhta  :)R=HRlM5#RsEHo0M_H8,CGRosHEH0_MG8C2R;R-O-RNE0OR0DHCDsN#R
RRNRPsLHNDsCRCD#k0RRRRRRRR:RRR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFIRV2=R:
RRRR5RRFC0Es=#R>jR''
2;RRRRPHNsNCLDRCXs#0kDRRRRRRRRRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRIRV-NoksL8_H20#R
:=RRRRRFR50sEC#>R=R''j2R;
RPRRNNsHLRDCb#sCkRD0RRRRRRRR: R)q
p;RCRLo
HMRRRR-Q-RVCRMoHN0PFCRskRMDsDRNCMo,CRs0Mks3R
RRVRHRC5DVH0_MG8CRV<RI02RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RHRRVNR5s<oRRjj32ER0CRM
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"mw_zQ7X :CRhoHN0PNCRslokCRM0b#N#C"8R
RRRRRRRR)&R 'qpHolNCs5No#2RCsPCHR0$CFsssR;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RRRRb#sCkRD0:N=Rs
o;RRRRHbVRskC#D>0R=.R53*j*5VDC0M_H8+CG4R220MEC
RRRRNRR#s#C0mRh_)WqhtQhRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"mw_zQ7X 5q) pR2:P0COF0sRsOkMN80C"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRVRHRCFPsFVDI0_#$RDC=HRVG_C8IbsNRC0EMR
RRRRRRsRbCD#k0=R:RCbs#0kDR8lFR35.j5**D0CV_8HMC4G+2R2;RR--IbsN
RRRRCRRD
#CRRRRRRRRskC0s#MRNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;
RRRRR8CMR;HV
RRRR8CMR;HV
RRRRsVFRHHRMsRXCD#k0N'sMRoCDbFF
RRRRHRRVsRbCD#k0=R>Rj.3*R*H0MEC
RRRRRRRRCXs#0kD5RH2:'=R4
';RRRRRRRRb#sCkRD0R:RR=sRbCD#k0RR-.*3j*
H;RRRRRDRC#RC
RRRRRXRRskC#DH052=R:R''j;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RRVRHRNoksL8_HR0#>RRjNRM8sMFk80_#$RDC=HRVG_C8sMFk8ER0CRM
RRRRR#sCkRD0:s=RF8kM_GVHC58RNRso=X>RskC#D50RD0CV_8HMCRG
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0sFRH0oE_8HMC,G2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCRslMNH8RCs=X>RskC#D50RsEHo0M_H8-CG4FR8IFM0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8-CGoskN8H_L0,#2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRR#CDCR
RRRRRskC#D:0R=sRXCD#k0sR5CD#k0N'sM2oC;R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0kF_VCHG8
;
RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRq) pR;RR-RR-CRsNRD
RORRF0M#NRM0D0CV_8HMCRGRR:RRRaQh )t ;-RR-CRDVH0RMG8CRH5EoHERMG8C2R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hat; )R-R-RosHEH0RMG8C
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C;RRRRO#FM00NMRNoksL8_HR0#RRRR:qRhaqz)pRRRRRRRRRRRRRRRRRRR:V=RH8GC_NoksL8_H20#R-R-RFyRVkRoNRs8L#H0
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0VRIRR:RRRaQh )t RR:=l#HMRH5so_E0HCM8Gs,RH0oE_8HMC;G2R-R-R0ONODERHs0CN
D#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0VFRI:2R=R
RRRRR5EF0CRs#='>Rj;'2
RRRRsPNHDNLCsRXCD#k0RR:z h)1emp #7_VCHG8DR5C_V0HCM8GR+48MFI0VFRIk-oN_s8L#H02=R:
RRRR5RRFC0Es=#R>jR''
2;RRRRPHNsNCLDRCbs#0kDR):R ;qp
LRRCMoH
RRRRRHV5VDC0M_H8RCG<IRV2ER0CRMRRRRRRRRRRR--MDkDRMsNoRC
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRVRHRs5No=R>R35.jD**C_V0HCM8GF2RssRNoRR<-35.jD**C_V0HCM8GR220MEC
RRRRNRR#s#C0mRh_)WqhtQhRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"mw_1Q7X 5q) pR2:P0COF0sRsOkMN80C"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRVRHRCFPsFVDI0_#$RDC=HRVG_C8#kN0sCN0RC0EMR
RRRRRRVRHRoNsRj<R30jRERCMRRRRRRRRRRRRR-R-R0#Nk0sNCR
RRRRRRRRRskC#D:0R=FRM0NR#0Nks05CRskC#DE0'H,oER#sCk'D0D2FI;RRRRRRRRR--kCM8sFVDIR
RRRRRRDRC#RC
RRRRRRRRR#sCkRD0:#=RNs0kNR0C5#sCk'D0EEHo,CRs#0kD'IDF2R;RRRRRRRRRR-R-RCFPsFVDIR
RRRRRRMRC8VRH;R
RRRRRRCRs0MksR#sCk;D0
RRRRCRRD
#CRRRRRRRRb#sCkRD0:N=RLN#5sRo2lRF85j.3*D*5C_V0HCM8G2+42R;RRRRRRRRRR-RR-sRINRb
RRRRR8CMR;HV
RRRR#CDCR
RRRRRb#sCkRD0:N=RLN#5s;o2
RRRR8CMR;HV
RRRRsVFRHHRMsRXCD#k0N'sMRoCDbFF
RRRRHRRVsRbCD#k0=R>Rj.3*R*H0MEC
RRRRRRRRCXs#0kD5RH2:'=R4
';RRRRRRRRb#sCkRD0R:RR=sRbCD#k0RR-.*3j*
H;RRRRRDRC#RC
RRRRRXRRskC#DH052=R:R''j;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RRVRHRoNsRj<R30jRE
CMRRRRRsRXCD#k0=R:R_0FVCHG805-F5_#X#sCk2D0,sRXCD#k0H'EoRE,X#sCk'D0D2FI;R
RRMRC8VRH;R
RRVRHRNoksL8_HR0#>RRjNRM8sMFk80_#$RDC=HRVG_C8sMFk8ER0CRM
RRRRR#sCkRD0:s=RF8kM_GVHC58RNRso=X>RskC#D50RD0CV_8HMCRG
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0sFRH0oE_8HMC,G2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCRslMNH8RCs=X>RskC#D50RsEHo0M_H8-CG4FR8IFM0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8-CGoskN8H_L0,#2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRR#CDCR
RRRRRskC#D:0R=sRXCD#k0sR5CD#k0N'sM2oC;R
RRMRC8VRH;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0#F_VCHG8
;
RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;RRRRRRRRRRRR-R-R#kMHCoM8R
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )R-R-RVDC0MRH8RCG5oEHEMRH82CG
RRRRMOF#M0N0HRso_E0HCM8GRRRRQ:Rhta  R)RRRRRRRRRRRRRRRRRRR:=jR;R-s-RH0oER8HMCRG
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMRtq)_wp aRR:Q hatR ):q=R)Dt'C0MoE;-4
RRRRHNDNX#RqR)tRRRRR:RRR)zh p1me_ 7zQh1t7h 5tq)_wp aFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDR#sCkRD0RRR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RoLCHRM
RHRRVsRNoC'DMEo0R4<RRRFs5VDC0M_H8RCG<HRso_E0HCM8G02RE
CMRRRRRCRs0MksRzhqwR;
RCRRMH8RVR;
RsRRCD#k0=R:R#sCHRxC5oNsRRRRRRRRRRRR=z>Rh1) m pe7V_kH8GCRq5X),t2
RRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=RVDC0M_H8,CG
RRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=RosHEH0_MG8C,R
RRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFR0_HkVG;C8
R
R-O-RFCMPs80CRsPC#MHF
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRso:hRz)m 1p7e _1zhQ th7R2RRRRRRRRR-k-RMo#HM
C8RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRFROMN#0Mq0R)pt_ Rwa:hRQa  t)=R:Rtq)'MDCo-0E4R;
RNRRD#HNR)XqtRRRRRRRRz:Rh1) m pe7h_z1hQt q75)pt_ Rwa8MFI0jFR2#RHRtq);R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR40MEC
RRRRsRRCs0kMqRhz
w;RRRRCRM8H
V;RRRRskC0szMRh1) m pe7V_kH8GC5sGNo
2;RMRC8kRVMHO0F0MRFV_kH8GC;R

RMVkOF0HMFR0_H#VGRC85R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;RRRRRRRRRRRRRRR--#MHoCR8
RORRF0M#NRM0D0CV_8HMCRGRR:RRRaQh )t ;-RR-CRDVH0RMG8CRH5EoHERMG8C2R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hatR )RRRRRRRRRRRRRRRRR=R:RRj;RR--sEHo0MRH8
CGRRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRMOF#M0N0)Rqt _pw:aRRaQh )t RR:=q')tDoCM04E-;R
RRDRNHRN#Xtq)RRRRRRRR:hRz)m 1p7e _t1Qh5 7q_)tpa wRI8FMR0FjH2R#)RqtR;
RPRRNNsHLRDCskC#DR0RRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR4F5sRD0CV_8HMC<GRRosHEH0_MG8C2ER0CRM
RRRRR0sCkRsMhwq1;R
RRMRC8VRH;R
RRCRs#0kDRR:=sHC#x5CRNRsoRRRRRRRRR=RR>hRz)m 1p7e _H#VGRC85)Xqt
2,RRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>D0CV_8HMC
G,RRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>sEHo0M_H8,CG
RRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D=CR>PRFCDsVF#I_0C$D2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0F#GVHC
8;
-RR-FROMsPC0RC8P#CsH
FMRkRVMHO0F0MRFV_#H8GCRR5
RNRRs:oRR)zh p1me_ 71hQt R72RRRRRRRRR-RR-HR#o8MC
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0q_)tpa wRQ:Rhta  :)R=)RqtC'DMEo0-
4;RRRRNNDH#qRX)RtRRRRRRRR:z h)1emp 17_Q th7)5qt _pw8aRF0IMF2RjRRH#q;)t
LRRCMoH
RRRRRHVN'soDoCM0<ERR04RE
CMRRRRRCRs0MksR1hqwR;
RCRRMH8RVR;
RsRRCs0kMhRz)m 1p7e _H#VG5C8GoNs2R;
R8CMRMVkOF0HMFR0_H#VG;C8
R
RVOkM0MHFR_0F#GVHC58RNRso:hRz)m 1p7e _HkVG2C8R0sCkRsMz h)1emp #7_VCHG8#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCRs5NoH'Eo4E+RI8FMR0FN'soD2FI;R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR40MEC
RRRRsRRCs0kMqRh1
w;RRRRCRM8H
V;RRRRskC#D50RN'soEEHoRI8FMR0FN'soD2FIRR:=z h)1emp #7_VCHG8D5OCPNMCNO5s2o2;R
RRCRs#0kDRs5NoH'Eo4E+2RRRRRRRRRRRR:RR=jR''R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0F#GVHC
8;
-RR-CRAO#NkCVRFRC0ERHVNsRD$ObFlDNHO0RC8#HHxMsoRk#DCRRHM0RECVCHG8FRbH
M0R-R-RObN	CNo#ER0CR#CVOkM0MHF#sRNCsRbF8PHC08RFFROl0bkCER0CCRs#0kDRMsNo
C#R-R-RN GlCbD:R
R-#-RHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-#-RHNoMDVRk.RR:kGVHC58RcFR8IFM0R2-.;R
R-#-RHNoMDVRk4Dlk0.kVRk:RVCHG8kR5VCHG8H_Eo5ERd-,Rd',R*R',c-,R.82RF0IMFR
R-R-RRRRRRRRRRRRRRRRRRRRRRRRRRkRRVCHG8F_DIdR5,dR-,*R''c,R,.R-2
2;R-R-R4kVl0kDkRV.<k=RV*4RR.kV;R
R-e-RN8DHRNOEs0NOC:s#R''+,-R''',R*R',',/'R''sRRFs'R)'5lsC2',RlF'RsvR''lR5F,82
-RR-4R''sR5CbOHsNFODR2,',q'R''NRL5N#R2,',h'R''MR#5-VCHG8R2
RMVkOF0HMVRkH8GC_oEHEDR5C_V0HCM8Gs,RH0oE_8HMCRGRRQ:Rhta  
);RRRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRRRRRRRRRRRRRRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8C.s,RH0oE_8HMCRG.:hRQa  t)RRR:j=R2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRROCN#RCFbsHN0FHMR#R
RRRRRIMECR''+|-R''>R=R0sCkRsMlHNGlRkl5VDC0M_H8,CGRVDC0M_H8.CG2RR+4R;
RRRRRCIEM*R''RRRR=RR>CRs0MksRVDC0M_H8RCG+CRDVH0_MG8C.RR+4R;
RRRRRCIEM/R''RRRR=RR>CRs0MksRVDC0M_H8RCG-HRso_E0HCM8G
.;RRRRRERIC'MR4R'RRRRR=s>RCs0kMsR-H0oE_8HMCRG;RRRRRRRRRRRRRRRRR-RR-CRsOsHbFDON
RRRRIRRERCM'|)''Rs'RR=>skC0slMRHRM#5VDC0M_H8,CGRVDC0M_H8.CG2R;R-"-Rs"Cl
RRRRIRRERCM'|v''Rl'RR=>skC0slMRHRM#5VDC0M_H8,CGRVDC0M_H8.CG2R;R-"-Rl"F8
RRRRIRRERCMFC0EsR#RRR=>skC0sDMRC_V0HCM8GR;R-w-RFNsRLN#RM88RCkVNDR0
RCRRMO8RN;#C
CRRMV8Rk0MOHRFMkGVHCE8_H;oE

RRRkRVMHO0FkMRVCHG8F_DIDR5C_V0HCM8Gs,RH0oE_8HMCRGRRQ:Rhta  
);RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRRRRRRRRRRRRRRRRRB:R]qq)B)a RR:=';X'
RRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMC,G.RosHEH0_MG8C.RR:Q hatR )R=R:R
j2RRRRskC0sQMRhta  H)R#R
RLHCoMR
RRNRO#FCRbNCs0MHFR
H#RRRRRERIC'MR+R'|'R-'=s>RCs0kMHRlM5#RsEHo0M_H8,CGRosHEH0_MG8C.
2;RRRRRERIC'MR*R'RRRRR=s>RCs0kMHRso_E0HCM8GRR+sEHo0M_H8.CG;R
RRRRRIMECR''/RRRRR>R=R0sCkRsMsEHo0M_H8RCG-CRDVH0_MG8C.RR-4R;
RRRRRCIEM4R''RRRR=RR>CRs0MksRC-DVH0_MG8CR4-R;RRRRRRRRRRRRRRRRRRR-s-RCbOHsNFODR
RRRRRIMECR'')|''sR>R=R0sCkRsMl#HMRH5so_E0HCM8Gs,RH0oE_8HMC2G.;-RR-sR"C
l"RRRRRERIC'MRv''|lR'R=s>RCs0kMHRlM5#RsEHo0M_H8,CGRosHEH0_MG8C.R2;RR--"8lF"R
RRRRRIMECREF0CRs#R>R=R0sCkRsMsEHo0M_H8;CGR-R-RsVFR#NLR8NMRV8CN0kD
RRRR8CMR#ONCR;
R8CMRMVkOF0HMVRkH8GC_IDF;R
R
VRRk0MOHRFM#GVHCE8_HRoE5VDC0M_H8,CGRosHEH0_MG8CR:RRRaQh )t ;R
RRRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMRRRRRRRRRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMC,G.RosHEH0_MG8C.RR:Q hatR )R=R:R
j2RRRRskC0sQMRhta  H)R#R
RLHCoMR
RRNRO#FCRbNCs0MHFR
H#RRRRRERIC'MR+R'|'R-'=s>RCs0kMNRlGkHllDR5C_V0HCM8GD,RC_V0HCM8GR.2+;R4
RRRRIRRERCM'R*'RRRRRR=>skC0sDMRC_V0HCM8GRR+D0CV_8HMCRG.+;R4
RRRRIRRERCM'R/'RRRRRR=>skC0sDMRC_V0HCM8GRR-sEHo0M_H8.CGR4+R;R
RRRRRIMECR''4RRRRR>R=R0sCkRsM-osHEH0_MG8CR4+R;RRRRRRRRRRRRRRRRR--sHCObOsFNRD
RRRRRCIEM)R''s|''=RR>CRs0MksRMlH#DR5C_V0HCM8GD,RC_V0HCM8G;.2R-R-RC"slR"
RRRRRCIEMvR''l|''=RR>CRs0MksRVDC0M_H8.CG;RRRRRRRRRRRRRRRRRRRR-R-RF"l8R"
RRRRRCIEMqR''N|''=RR>CRs0MksRVDC0M_H8RCG+;R4RRRRRRRRRRRRRRRRR-R-RL"N#R"
RRRRRCIEMhR''M|''=RR>CRs0MksRVDC0M_H8RCG+;R4RRRRRRRRRRRRRRRRR-R-RV-#H8GC
RRRRIRRERCMFC0EsR#RRR=>skC0sDMRC_V0HCM8GR;
RCRRMO8RN;#C
CRRMV8Rk0MOHRFM#GVHCE8_H;oE
R
RVOkM0MHFRH#VG_C8DRFI5VDC0M_H8,CGRosHEH0_MG8CR:RRRaQh )t ;R
RRRRRRRRRRRRRRRRRRRRRRCFbsHN0FRMRRRRRRRRRRRRRR:RRRqB])aqB :)R=XR''R;
RRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8C.s,RH0oE_8HMCRG.:hRQa  t)RRR:j=R2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRROCN#RCFbsHN0FHMR#R
RRRRRIMECR''+|-R''>R=R0sCkRsMl#HMRH5so_E0HCM8Gs,RH0oE_8HMC2G.;R
RRRRRIMECR''*RRRRR>R=R0sCkRsMsEHo0M_H8RCG+HRso_E0HCM8G
.;RRRRRERIC'MR/R'RRRRR=s>RCs0kMHRso_E0HCM8GRR-D0CV_8HMC;G.
RRRRIRRERCM'R4'RRRRRR=>skC0s-MRD0CV_8HMCRG;RR--sHCObOsFNRD
RRRRRCIEM)R''s|''=RR>CRs0MksRMlH#sR5H0oE_8HMCRG,sEHo0M_H8.CG2R;R-"-Rs"Cl
RRRRIRRERCM'|v''Rl'RR=>skC0slMRHRM#5osHEH0_MG8C,HRso_E0HCM8G;.2R-R-RF"l8R"
RRRRRCIEM0RFE#CsR=RR>CRs0MksRosHEH0_MG8C;-RR-CR8VDNk0FRVsLRN#M,RCNoRM88RCkVNDR0
RCRRMO8RN;#C
CRRMV8Rk0MOHRFM#GVHCD8_F
I;
-RR-NR1lNCR#LRNF,PCR0LkRHk#M0oRE"CR#CHx_#sC"MRHbRk0F$MDRsVFRC0EHssRNCMo#R:
RR--#MHoNkDRVk4lDV0k.RR:kGVHC58RkGVHCE8_HRoE54kV,*R''k,RVR.28MFI0RF
RR--RRRRRRRRRRRRRRRRRRRRRRRRRRRRkGVHCD8_F5IRk,V4R''*,VRk.;22
-RR-VRk4Dlk0.kVRR<=kRV4*VRk.R;R
VRRk0MOHRFMkGVHCE8_HRoE5x#HCC_s#:RRR)zh p1me_ 7kGVHC
8;RRRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRR:B)]qq Ba)=R:R''X;R
RRRRRRRRRRRRRRRRRRRRRRHR#xsC_CR#.:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RsRRCs0kMVRkH8GC_oEHEDR5C_V0HCM8GRRR=#>RH_xCs'C#EEHo,R
RRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8G=RR>HR#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRR=>FsbCNF0HMR,
RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GR.R=#>RH_xCs.C#'oEHER,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRG.=#>RH_xCs.C#'IDF2R;
R8CMRMVkOF0HMVRkH8GC_oEHE
;
RkRVMHO0FkMRVCHG8F_DI#R5H_xCsRC#Rz:Rh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRRRRRRCFbsHN0F:MRRqB])aqB :)R=XR''R;
RRRRRRRRRRRRRRRRRRRRRHR#xsC_CR#.:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RsRRCs0kMVRkH8GC_IDFRC5DVH0_MG8CR=RR>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGRR=>#CHx_#sC'IDF,R
RRRRRRRRRRRRRRRRRRRRRRCFbsHN0FRMRR>R=RCFbsHN0F
M,RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GR.R=#>RH_xCs.C#'oEHER,
RRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8G=.R>HR#xsC_C'#.D2FI;R
RCRM8VOkM0MHFRHkVG_C8D;FI
R
RVOkM0MHFRH#VG_C8EEHoRH5#xsC_CR#R:hRz)m 1p7e _H#VG;C8
RRRRRRRRRRRRRRRRRRRRRRRRCFbsHN0F:MRRqB])aqB :)R=XR''R;
RRRRRRRRRRRRRRRRRRRRR#RRH_xCs.C#Rz:Rh1) m pe7V_#H8GC2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRRskC0s#MRVCHG8H_Eo5ERD0CV_8HMCRGRRR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGR=#>RH_xCs'C#D,FI
RRRRRRRRRRRRRRRRRRRRRRRRCFbsHN0FRMRR>R=RCFbsHN0F
M,RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRG.RR=>#CHx_#sC.H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8.CGRR=>#CHx_#sC.F'DI
2;RMRC8kRVMHO0F#MRVCHG8H_Eo
E;
VRRk0MOHRFM#GVHCD8_F5IR#CHx_#sCRRR:z h)1emp #7_VCHG8R;
RRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFM:]RBqB)qaR ):'=RX
';RRRRRRRRRRRRRRRRRRRRR#RRH_xCs.C#Rz:Rh1) m pe7V_#H8GC2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRRskC0s#MRVCHG8F_DIDR5C_V0HCM8GRRR=#>RH_xCs'C#EEHo,R
RRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CR>R=Rx#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRbRFC0sNHRFMR=RR>bRFC0sNH,FM
RRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRG.RR=>#CHx_#sC.H'Eo
E,RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRG.=#>RH_xCs.C#'IDF2R;
R8CMRMVkOF0HMVR#H8GC_IDF;R

RR--bbksF:#CR0sCk#sMR#NRNs0kN80CRlMkL
CsRkRVMHO0F#MRNs0kNR0C5R
RRFROMN#0MD0RC_V0HCM8G:RRRaQh )t ;R
RRFROMN#0Ms0RH0oE_8HMC:GRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMR0#NRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CGR
:=RRRRRFR50sEC#>R=R''42R;
RoLCHRM
RsRRCs0kMNR#0R;
R8CMRMVkOF0HMNR#0Nks0
C;
-RR-kRbs#bFCs:RCs0kMN#RR0#Nk0sNCM8RkClLsR
RVOkM0MHFR0#Nk0sNC
R5RRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHND#CRN:0RR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G:2R=R
RRRRR5EF0CRs#='>R4;'2
LRRCMoH
RRRRR--#kN0sCN0R#bFHP0HC0,RFNR#0Nks0MCRC0oNH,PCR#[k0FR8RF"M0NR#0Nks02C5"R
RRNR#0DR5C_V0HCM8G:2R=jR''R;
RsRRCs0kMNR#0R;
R8CMRMVkOF0HMNR#0Nks0
C;
VRRk0MOHRFM#kN0sCN0RR5
R#RRH_xCsRC#:hRz)m 1p7e _HkVG2C8RRRRR-RR-MRFD0$RE#CRHRxCF0VRERH#Hk#R#
C8RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s#MRNs0kNR0C5x#HCC_s#H'EoRE,#CHx_#sC'IDF2R;
R8CMRMVkOF0HMNR#0Nks0
C;
VRRk0MOHRFM#kN0sCN0RR5
R#RRH_xCsRC#:hRz)m 1p7e _H#VG2C8RRRRR-RR-MRFD0$RE#CRHRxCF0VRERH#Hk#R#
C8RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s#MRNs0kNR0C5x#HCC_s#H'EoRE,#CHx_#sC'IDF2R;
R8CMRMVkOF0HMNR#0Nks0
C;
-RR-#RqRONRFCMO#F#HMFR0RF0E#ICREkFR#NCRRNosbOEHN7DR1CuRMsPHFCMlM
0,R-R-RC0E#VCRk0MOH#FMR	0NCNRbsCNl0#CsRRHM0#EFCFR0FRD#VlFsNN0RMO8Rs0CNCR
R-V-RH8GCRHbFMM0RkClLsR#3RCaE#VCRk0MOH#FMRCNsR#8CHCoM8FR0RMOFP0CsRFVslR
R-N-RR8#0_oDFHPO_CFO0sFR0RC0ER7e]pHRVGRC8bMFH0FRVs0lNRHk#M0oREOCRFCMPMF0HMR#
RR--F0VRECC#RObN	CNo#R3RQNMRRsbkC]Re7CpRMsPHFCMlM$0RF#kREDFk8#RkCER0CR
R-"-R0kF_VCHG8N"RM"8R0#F_VCHG8s"RFHk0M3C#
-RR-MRz#MHoCV8RH8GCRHbFMR0
RMVkOF0HMFR0_HzwG
R5RRRRNRsoRRRRR1:Raz7_pQmtB _eB)am;R
RRHRI8R0ER:RRRahqzp)q;RRRRRRRRRRRRRRRR-R-R8IH0FERVCRPOs0F
RRRRNVsOF0HMRR:hzqa)2qpRRRRRRRRRRRRRRRRRR--I0H8EVRFRNVsOF0HMR
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC858IH0VE-s0NOH-FM4FR8IFM0Rs-VNHO0F;M2
LRRCMoH
RRRRRHV5oNs'MDCoR0E/s=RCD#k0C'DMEo02ER0CRM
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"mw_zQ5XR1_a7ztpmQeB_ mBa)"2R
RRRRRRRR"&Re0COFDsRC0MoE8#RFFRM0NRl03OERMRQbRk0DoCM0HER#
R"RRRRRRRR&hRQa  t)l'HN5oCN'soDoCM0RE2&RR"NRM8Fbk0kI0RHRDDL"CR
RRRRRRRRQ&Rhta  H)'lCNo5#sCk'D0DoCM0RE2&RR"ICH83R"
RRRRR#RRCsPCHR0$CFsssR;
RRRRR0sCkRsMhwqz;R
RRDRC#RC
RRRRR#sCkRD0:0=RFV_kH8GCRs5Nos,RCD#k0H'EoRE,skC#DD0'F;I2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FzGwH;R

RR--#MHoCV8RH8GCRHbFMR0
RMVkOF0HMFR0_H1wG
R5RRRRNRsoRRRRR1:Raz7_pQmtB _eB)am;R
RRHRI8R0ER:RRRahqzp)q;RRRRRRRRRRRRRRRR-R-R8IH0FERVCRPOs0F
RRRRNVsOF0HMRR:hzqa)2qpRRRRRRRRRRRRRRRRRR--I0H8EVRFRNVsOF0HMR
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC858IH0VE-s0NOH-FM4FR8IFM0Rs-VNHO0F;M2
LRRCMoH
RRRRRHV5oNs'MDCoR0E/s=RCD#k0C'DMEo02ER0CRM
RRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"mw_1Q5XR1_a7ztpmQeB_ mBa)"2R
RRRRRRRR"&Re0COFDsRC0MoE8#RFFRM0NRl03OERMRQbRk0DoCM0HER#
R"RRRRRRRR&hRQa  t)l'HN5oCN'soDoCM0RE2&RR"NRM8Fbk0kI0RHRDDL"CR
RRRRRRRRQ&Rhta  H)'lCNo5#sCk'D0DoCM0RE2&RR"ICH83R"
RRRRR#RRCsPCHR0$CFsssR;
RRRRR0sCkRsMhwq1;R
RRDRC#RC
RRRRR#sCkRD0:0=RFV_#H8GCRs5Nos,RCD#k0H'EoRE,skC#DD0'F;I2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0F1GwH;R

RR--V8HMHRMo0RECLMFk8F#RVRRNMLklCRs3RCaE#VCRk0MOH#FMRMONRRLCk8#CR	DHCER0H
#:R-R-Ro#HMRNDGRGG:VRkH8GCRR5(8MFI0-FRd
2;R-R-RR--WOEHE#RHRC0ERl#NC#RNRV"kH8GCRw5zHEG_HRoE5,44d82RF0IMFwRzHDG_F4I542,d2R"
RR--#MHoN$DR$:$RRHkVGRC85HzwGH_Eo5ER4R4,d",R+R",4R4,dR2
RR--RRRRRRRRRRRRRFR8IFM0RHzwGF_DI454,,RdR""+,4R4,2Rd2R;
RR--WsECC4R"4H"R#ER0CHRI8R0EFGVRG5GRG'GGDoCM0,E2
-RR-MRN8RRdH0#REDCRFsICRkLFM58RNRL#5GGG'IDF2R2
RR--QNMRRsbkC]Re7CpRMsPHFCMlMk0R#"CRkGVHCE8_H"oER8NMRV"kH8GC_IDF"R
RVOkM0MHFRHkVGH_Eo5ER
RRRR8IH0RE,VOsN0MHFR:RRRahqzp)q;R
RRbRFC0sNHRFMRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRI0H8ER.,VOsN0MHF.RR:hzqa)RqpR=R:R
j2RRRRskC0sQMRhta  H)R#R
RLHCoMR
RRCRs0MksRHkVG_C8EEHoRC5DVH0_MG8CR=RR>HRI8R0E-RR4-sRVNHO0F
M,RRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGRR=>-NVsOF0HMR,
RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRRRR=F>RbNCs0MHF,R
RRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8C.=RR>HRI8.0ER4-RRV-Rs0NOH.FM,R
RRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8G=.R>VR-s0NOH.FM2R;
R8CMRMVkOF0HMVRkHEG_H;oE
R
RVOkM0MHFRHkVGF_DI
R5RRRRI0H8EV,Rs0NOHRFMRRR:hzqa);qp
RRRRCFbsHN0FRMRRRRRR:RRRqB])aqB :)R=XR''R;
RIRRHE80.V,Rs0NOH.FMRh:Rq)azqRpRRR:=jR2
RsRRCs0kMhRQa  t)#RH
LRRCMoH
RRRR0sCkRsMkGVHCD8_F5IRD0CV_8HMCRGRRR=>I0H8ERR-4RR-VOsN0MHF,R
RRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CR>R=Rs-VNHO0F
M,RRRRRRRRRRRRRRRRRRRRRFRRbNCs0MHFRRRR=F>RbNCs0MHF,R
RRRRRRRRRRRRRRRRRRRRRRVDC0M_H8.CGR>R=R8IH0RE.-RR4-sRVNHO0F,M.
RRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8.CGRR=>-NVsOF0HM;.2
CRRMV8Rk0MOHRFMkGVH_IDF;R

RMVkOF0HMVR#HEG_HRoE5R
RRHRI8,0ERNVsOF0HMRRR:qRhaqz)pR;
RFRRbNCs0MHFRRRRRRRRRB:R]qq)B)a RR:=';X'
RRRR8IH0,E.RNVsOF0HM:.RRahqzp)qR:RR=2Rj
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RsRRCs0kMVR#H8GC_oEHEDR5C_V0HCM8GRRR=I>RHE80RV-Rs0NOH,FM
RRRRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CR>R=Rs-VNHO0F
M,RRRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRR=>FsbCNF0HMR,
RRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GR.R=I>RHE80.RR-VOsN0MHF.R,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRG.=->RVOsN0MHF.
2;RMRC8kRVMHO0F#MRV_HGEEHo;R

RMVkOF0HMVR#HDG_F5IR
RRRR8IH0RE,VOsN0MHFR:RRRahqzp)q;R
RRbRFC0sNHRFMRRRRRRRR:]RBqB)qaR ):'=RX
';RRRRI0H8ER.,VOsN0MHF.RR:hzqa)RqpR=R:R
j2RRRRskC0sQMRhta  H)R#R
RLHCoMR
RRCRs0MksRH#VG_C8DRFI5VDC0M_H8RCGR>R=R8IH0-ERRNVsOF0HMR,
RRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8G=RR>VR-s0NOH,FM
RRRRRRRRRRRRRRRRRRRRRRRFsbCNF0HMRRRRR=>FsbCNF0HMR,
RRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8C.=RR>HRI8.0ERV-Rs0NOH.FM,R
RRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8C.>R=Rs-VNHO0F2M.;R
RCRM8VOkM0MHFRH#VGF_DI
;
RkRVMHO0F0MRFM_k#MHoC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-VRkH8GCRHbFMH0RM0bk
RRRRMOF#M0N0HR#xRCRRRRRRRRRRh:Rq)azqRp;RRRRRRRRR-RR-CRDMEo0RRFVFbk0kR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0s0MRFM_k#C5s#CHxRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=Rx#HC,-4
RRRRRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=R
j,RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRFRRPVCsD_FI#D0$C>R=RCFPsFVDI0_#$2DC2R;
R8CMRMVkOF0HMFR0_#kMHCoM8
;
RkRVMHO0F0MRFM_k#MHoC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;RRRRR--kGVHCb8RF0HMRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;-RR-CRDMEo0RRFVFbk0kR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0s0MRFM_k#MHoC58RNRsoRRRRRRRRR=RR>sRNoR,
RRRRRRRRRRRRRRRRRRRRR#RRHRxCRRRRRRRRR>R=Rx#HCC_s#C'DMEo0,R
RRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RMRC8kRVMHO0F0MRFM_k#MHoC
8;
VRRk0MOHRFM0#F_HCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RH#VGRC8bMFH0MRHb
k0RRRRO#FM00NMRx#HCRRRRRRRRRRR:qRhaqz)pR;RRRRRRRRRR-R-RMDCoR0EFFVRkk0b0R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$2DC
RRRR0sCkRsMz h)1emp 17_Q th7#RH
LRRCMoH
RRRR0sCkRsM0#F_5#sCHRxC5oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>HR#x4C-,R
RRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>jR,
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D2C2;R
RCRM8VOkM0MHFR_0F#MHoC
8;
VRRk0MOHRFM0#F_HCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8R-R-RH#VGRC8bMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh; 7R-R-RCk#8FRVsCRDMEo0RRFVFbk0kR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR_0F#MHoC58RNRsoRRRRRRRRR=RR>sRNoR,
RRRRRRRRRRRRRRRRRRRRRx#HCRRRRRRRRRRR=#>RH_xCs'C#DoCM0
E,RRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRFRRPVCsD_FI#D0$C>R=RCFPsFVDI0_#$2DC;R
RCRM8VOkM0MHFR_0F#MHoC
8;RRR
RMVkOF0HMFR0_NsCD
R5RRRRNRso:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRR-k-RVCHG8FRbHRM0HkMb0R
RRCRs0MksRq) pR
RHR#
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)=R:RoNs'oEHER;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)=R:RoNs'IDF;R
RRNRPsLHNDsCRCD#k0RRRR:RRRq) pR;RRRRRR-R-R#sCk
D0RRRRPHNsNCLDRoNs_0HMRRRRRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RLHCoMR
RRVRHRs5NoC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMj;3j
RRRR8CMR;HV
RRRRoNs_0HMRR:=0GF_jO45DMCNP5CON2so2R;
RHRRVQR5#5_XN_soH2M02ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"_am)p qRV5kH8GC2l:RCP0NNCDkR08CCCO08s,RCs0kMoHMRjj3"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRjj3;R
RRMRC8VRH;R
RRCRs#0kDRR:=j;3j
RRRRsVFRHHRMsRNoM_H0N'sMRoCDbFF
RRRRHRRVNR5sHo_MH052RR='24'RC0EMR
RRRRRRCRs#0kDRR:=skC#D+0RR35.jH**2R;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FsDCN;R

RMVkOF0HMFR0_NsCD
R5RRRRNRso:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRR-k-RVCHG8FRbHRM0HkMb0R
RRCRs0MksRq) pR
RHR#
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)=R:RoNs'oEHER;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)=R:RoNs'IDF;R
RRNRPsLHNDsCRCD#k0RRRR:RRRq) pR;RRRRRR-R-R#sCk
D0RRRRPHNsNCLDRoNs_0HMRRRRRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RR-R-R#kMHCoM8CRPsF#HMVRFRoNskMlC0R
RRNRPsLHNDNCRsko_MR#RR:RRR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRR-N-RLD#FkR0CFNVRslokC
M0RCRLo
HMRRRRH5VRN'soDoCM0<ERRR420MEC
RRRRsRRCs0kM3RjjR;
RCRRMH8RVR;
RNRRsHo_M:0R=FR0_4Gj5CODNCMPOs5No;22
RRRRRHV5_Q#Xs5NoM_H0R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"m _)q5pR#GVHC:82R0lCNDPNk8CRCO0C0,C8R0sCkHsMMjoR3
j"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sjMR3
j;RRRRCRM8H
V;RRRRN_sokRM#:0=RFV_kH8GCRs5NoM_H0
2;RRRRskC#DR0R:0=RFC_sN5DRN_sok2M#;R
RRVRHRs5NoM_H0s5NoM_H0H'EoRE2=4R''02RE
CMRRRRRCRs#0kDRR:=-#sCk;D0
RRRR8CMR;HV
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F0MRFC_sN
D;
VRRk0MOHRFM0HF_Mo0CC5sR
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_kH8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMqRhaqz)pR
RHR#
RORRF0M#NRM0D0CV_8HMC:GRRaQh )t RR:=N'soEEHo;R
RRNRPsLHNDNCRsko_MR#RRRR:z h)1emp z7_ht1QhR 75VDC0M_H8+CG4FR8IFM0R
j2RRRRR=R:R05FE#CsRR=>'2j';R
RLHCoMR
RRVRHRs5NoC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMjR;
RCRRMH8RVR;
RHRRVQR5#R_X5oNs202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR&RRRm"a_aQh )t RV5kH8GC2l:RCP0NNCDkR08CCCO08s,RCs0kMoHMR
j"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0sjMR;R
RRMRC8VRH;R
RRVRHRC5DVH0_MG8CR-<R402RE
CMRRRRRCRs0MksR
j;RRRRCRM8H
V;RRRRN_sokRM#:0=RFM_k#C5s#CHxRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=RoNs_#kM'oEHER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CRRRR=j>R,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C;22
RRRR0sCkRsM0HF_Mo0CC5sRN_sok2M#;R
RCRM8VOkM0MHFR_0FHCM0o;Cs
R
RVOkM0MHFR_0FHCM0oRCs5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-V-RH8GCRHbFMH0RM0bk
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0sQMRhta  R)
R
H#RRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  :)R=sRNoH'Eo
E;RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  :)R=sRNoF'DIR;
RPRRNNsHLRDCN_so#RRRRRRR:hRz)m 1p7e _t1QhR 75VDC0M_H8+CG4FR8IFM0R;j2
LRRCMoH
RRRRRHV5oNs'MDCoR0E<2R4RC0EMR
RRRRRskC0sjMR;R
RRMRC8VRH;R
RRVRHR#5Q_5XRN2so2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"_amQ hatR )5H#VG2C8:CRl0NNPDRkC8CC0O80C,CRs0MksHRMojR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kM;Rj
RRRR8CMR;HV
RRRRRHV5VDC0M_H8RCG<4R-2ER0CRM
RRRRR0sCkRsMjR;
RCRRMH8RVR;
RNRRs#o_RR:=0#F_5#sCHRxC5oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>N_so#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>jR,
RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D2C2;R
RRCRs0MksR_0FHCM0oRCs5oNs_;#2
CRRMV8Rk0MOHRFM0HF_Mo0CC
s;
VRRk0MOHRFM0jF_4
R5RRRR#RRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;RRRRRRRRRRRRR-k-RVCHG8FRbHRM0HkMb0R
RRFROMN#0MX0RvRqu:aR17p_zmBtQRR:='2j'RRRRRRRRRRRRR-R-RbvNR0GRFR
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85s#'NCMo2R;R-s-RCD#k0R
RLHCoMR
RRVRHR'5#DoCM0<ERRR420MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRR&aR"m4_j5HkVG2C8:kRMD8DRCO0C0,C8R0sCkHsMMhoRz"pp
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMhwqz;R
RRMRC8VRH;R
RRCRs0MksR_0FVCHG80R5F4_j5_0Fk5M##R2,Xuvq2#,R'oEHE#,R'IDF2R;
R8CMRMVkOF0HMFR0_;j4
R
RVOkM0MHFR_0Fj54R
RRRRR#RRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--#GVHCb8RF0HMRbHMkR0
RORRF0M#NRM0XuvqR1:Raz7_pQmtB=R:R''j2-RR-NRvbRRG0RF
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCR'5#soNMC
2;RCRLo
HMRRRRH5VR#C'DMEo0R4<R2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRR&"_amj#45VCHG8R2:MDkDR08CCCO08s,RCs0kMoHMRphzpR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMqRh1
w;RRRRCRM8H
V;RRRRskC0s0MRFH_VGRC85_0Fj045F5_##R2,Xuvq2#,R'oEHE#,R'IDF2R;
R8CMRMVkOF0HMFR0_;j4
R
RVOkM0MHFR_Q#X
R5RRRRNRso:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMApmm 
qhR#RH
RRRRsPNHDNLCsRNoP#DR1:Raz7_pQmtB _eB)amRs5NoC'DMEo0-84RF0IMF2Rj;-RR-DR#PR
RLHCoMR
RRsRNoP#DRR:=0#F_k5DPN2so;R
RRCRs0MksR_Q#XNR5sDo#P
2;RMRC8kRVMHO0FQMR#;_X

RRRkRVMHO0FQMR#R_X5R
RRsRNoRR:z h)1emp #7_VCHG8R2
RsRRCs0kMmRAmqp hR
RHR#
RPRRNNsHLRDCN#soD:PRR71a_mzpt_QBea Bm5)RN'soDoCM04E-RI8FMR0FjR2;RR--#
DPRCRLo
HMRRRRN#soD:PR=FR0_D#kPs5No
2;RRRRskC0sQMR#R_X5oNs#2DP;R
RCRM8VOkM0MHFR_Q#X
;
RkRVMHO0FaMRFj_X4
R5RRRRNRso:hRz)m 1p7e _HkVG2C8
RRRR0sCkRsMz h)1emp k7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM0kF_VCHG8aR5Fj_X4F50_D#kPs5No,22RoNs'oEHEN,RsDo'F;I2
CRRMV8Rk0MOHRFMaXF_j
4;
VRRk0MOHRFM0XF_j54R
RRRRoNsRz:Rh1) m pe7V_#H8GC2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksR_0F#GVHC58RaXF_j045Fk_#DNP5s2o2,sRNoH'EoRE,N'soD2FI;R
RCRM8VOkM0MHFR_aFX;j4
R
RVOkM0MHFR_aFXZj4RR5
RNRRs:oRR)zh p1me_ 7kGVHC
82RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s0MRFV_kH8GCRF5a_4XjZF50_D#kPs5No,22RoNs'oEHEN,RsDo'F;I2
CRRMV8Rk0MOHRFMaXF_j;4Z
R
RVOkM0MHFR_0FXZj4RR5
RNRRs:oRR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s0MRFV_#H8GCRF5a_4XjZF50_D#kPs5No,22RoNs'oEHEN,RsDo'F;I2
CRRMV8Rk0MOHRFMaXF_j;4Z
R
RVOkM0MHFR_aFz4XjRR5
RNRRs:oRR)zh p1me_ 7kGVHC
82RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s0MRFV_kH8GCRF5a_jzX4F50_D#kPs5No,22RoNs'oEHEN,RsDo'F;I2
CRRMV8Rk0MOHRFMazF_X;j4
R
RVOkM0MHFR_0Fz4XjRR5
RNRRs:oRR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s0MRFV_#H8GCRF5a_jzX4F50_D#kPs5No,22RoNs'oEHEN,RsDo'F;I2
CRRMV8Rk0MOHRFMazF_X;j4

RRRkRVMHO0FsMRCx#HC
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8RRRRRRRRRRRR-H-RM0bk
RRRRMOF#M0N0CRDVH0_MG8CRRRRRQ:Rhta  R);RR--HCM0oRCsb0FsH
FMRRRRO#FM00NMRosHEH0_MG8CRRRR:hRQa  t)R;R-#-RHRxCFVVRs0NOH
FMRRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRMOF#M0N0sRNooEHERR:Q hatR ):l=RNlGHk5lRN'soEEHo,sRNoF'DI
2;RRRRO#FM00NMRoNsDRFIRQ:Rhta  :)R=HRlM5CRN'soEEHo,sRNoF'DI
2;RRRRPHNsNCLDRPHMCRORRz:Rh1) m pe7V_kH8GCRs5NooEHEFR8IFM0RoNsD2FI;R
RRNRPsLHNDsCRCD#k0:RRR)zh p1me_ 7kGVHCD85C_V0HCM8GFR8IFM0RosHEH0_MG8C2=R:
RRRR5RRFC0Es=#R>jR''
2;RRRRPHNsNCLDRCMC8s#_F8kMHRMo:mRAmqp h=R:RDVN#
C;RCRLoRHMRR--sHC#xRC
RHRRVNR5sDo'C0MoERR<4F2RssR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwqz;R
RRDRC#RHV5PHMCDO'C0MoERR<402RE
CMRRRRRCRs0MksR#sCk;D0RRRRRRRRRRRRRRRRRRRR-#-R0MsHoHRD0NCsDNRPD
kCRRRRCCD#
RRRRHRRMOPCRR:=ONDCMOPC5oNs2R;
RRRRRRHV5osHEH0_MG8CRN>RsHoEoRE20MECR-RR-CRs0MksRb0FRsxCFR#
RRRRRMRRC#C8_ksFMM8Ho=R:RF5sk_M8#D0$CRR=VCHG8F_sk2M8R8NM
RRRRRRRRRRRRRRRRRRRRRRRR5RRsEHo0M_H8RCG=sRNooEHE2+4;R
RRRRRCHD#VDR5C_V0HCM8GRR<NDsoFRI20MECR-R-R0sCkRsMFsPCVIDF
RRRRRRRRRHV5CFPsFVDI0_#$RDC=HRVG_C8#kN0sCN02MRN8R
RRRRRRRRR55Fs0#F_k5DPHCMPOR22=4R''02RE
CMRRRRRRRRRCRs#0kDRR:=#kN0sCN0RC5s#0kD'oEHEs,RCD#k0F'DIR2;RRRR-#-RNs0kN
0CRRRRRRRRCRM8H
V;RRRRRDRC#RHV5oNsEEHoRD>RC_V0HCM8G02RE
CMRRRRRRRR-I-RsRNbF#sRNs0kN?0C
RRRRRRRRRHV5CFPsFVDI0_#$RDC=HRVG_C8#kN0sCN0R8NM
RRRRRRRRRRRRRFs5_0F#PkD5PHMCNO5sHoEo8ERF0IMFCRDVH0_MG8C+2422RR='24'
RRRRRRRRC0EMR
RRRRRRRRRskC#D:0R=NR#0Nks05CRskC#DE0'H,oER#sCk'D0D2FI;RRRR-R-R0#Nk0sNCR
RRRRRRDRC#RC
RRRRRRRRRRHV5oNsDRFI>s=RH0oE_8HMCRG20MEC
RRRRRRRRRRRR#sCkRD05VDC0M_H8RCG8MFI0NFRsFoDI:2R=R
RRRRRRRRRRRRRHCMPOC5DVH0_MG8CRI8FMR0FNDsoF;I2
RRRRRRRRCRRD
#CRRRRRRRRRRRRskC#D50RD0CV_8HMC8GRF0IMFHRso_E0HCM8G:2R=R
RRRRRRRRRRRRRHCMPODR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RRRRRRRRRMRRC#C8_ksFMM8Ho=R:RF5sk_M8#D0$CRR=VCHG8F_sk2M8;-RR-FRsk
M8RRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R
RRRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RoNsEEHoRR<=HCM0oRCsI0H8ER
RRRRRRVRHRs5NoIDFRR>=sEHo0M_H82CGRC0EMR
RRRRRRRRRskC#D50RNEsoHRoE8MFI0NFRsFoDI:2R=MRHP;CO
RRRRRRRR#CDCR
RRRRRRRRRskC#D50RNEsoHRoE8MFI0sFRH0oE_8HMCRG2:R=
RRRRRRRRRHRRMOPCRs5NooEHEFR8IFM0RosHEH0_MG8C2R;
RRRRRRRRRCMC8s#_F8kMHRMo:5=RsMFk80_#$RDC=HRVG_C8sMFk8R2;R-RR-FRsk
M8RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRRRR-)-RF8kMR#sCk
D0RRRRRVRHRCMC8s#_F8kMHRMo0MEC
RRRRRRRR#sCkRD0:s=RF8kM_GVHC58RNRsoRRRRRRRRR=RR>CRs#0kD,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlsCN8HMCRsRRRRR=H>RMOPCRH5so_E0HCM8G
-4RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0NFRsFoDI
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRRPVCsD_FI#D0$C>R=RCFPsFVDI0_#$2DC;R
RRRRRCRM8H
V;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFMsHC#x
C;
VRRk0MOHRFMsHC#x5CR
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_#H8GC;RRRRRRRR-RR-MRHb
k0RRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-H-RMo0CCbsRFHs0FRM
RORRF0M#NRM0sEHo0M_H8RCGR:RRRaQh )t ;-RR-HR#xFCRVsRVNHO0FRM
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0D
C;RRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D2R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRO#FM00NMRoNsEEHoRQ:Rhta  :)R=NRlGkHllNR5sEo'H,oERoNs'IDF2R;
RORRF0M#NRM0NDsoFRIR:hRQa  t)=R:RMlHCNR5sEo'H,oERoNs'IDF2R;
RPRRNNsHLRDCHCMPORRR:hRz)m 1p7e _H#VGRC85oNsEEHoRI8FMR0FNDsoF;I2
RRRRsPNHDNLCCRs#0kDRRR:z h)1emp #7_VCHG8C5DVH0_MG8CRI8FMR0FsEHo0M_H82CGR
:=RRRRRFR50sEC#>R=R''j2R;
RPRRNNsHLRDCskC8ORC8RRRRR:RRR71a_mzpt;QB
RRRRsPNHDNLCCRMC_8#sMFk8oHMRA:Rm mpq:hR=NRVD;#CRRRRRRRRR-RR-FRskHM8MRo
RoLCHRMR-s-RCx#HCR
RRVRHRs5NoC'DMEo0R4<R2sRFRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;1w
RRRR#CDH5VRHCMPOC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMskC#DR0;RRRRRRRRRRRRRRRRR-RR-0R#soHMR0DHCDsNRDPNkRC
RCRRD
#CRRRRRMRHPRCO:O=RDMCNP5CON2so;R
RRRRRH5VRsEHo0M_H8RCG>sRNooEHE02RERCMR-R-R0sCkRsM0RFbxFCs#R
RRRRRRVRHRs5NoF'DI=R/RaQh )t 'IDF2ER0CRMR-O-RE	CORsVFRDNRHs0CNRD
RRRRRRRRR#sCkRD0:5=RFC0Es=#R>sRNos5NooEHE;22RRRRRRRRRRRRRR--#MHoR0CGC
M8RRRRRRRRCRM8H
V;RRRRRRRRM8CC#F_skHM8M:oR=sR5F8kM_$#0D=CRRGVHCs8_F8kM2MRN8R
RRRRRRRRRRRRRRRRRRRRRRRRR5osHEH0_MG8CRN=RsHoEo4E+2R;
RRRRR#CDH5VRD0CV_8HMC<GRRoNsD2FIRC0EM-RR-CRs0MksRCFPsFVDIR
RRRRRRVRHRP5FCDsVF#I_0C$DRV=RH8GC_0#Nk0sNC02RE
CMRRRRRRRRRCRs8CkO8=R:RRFs5_0F#PkD5PHMC2O2;R
RRRRRRRRRH5VRskC8ORC8=4R''02RE
CMRRRRRRRRRRRRH5VRHCMPOs5NooEHE=2RR''j2ER0CRM
RRRRRRRRRRRRRR--#kN0sCN0R1umQeaQ R
RRRRRRRRRRRRRskC#D:0R=NR#0Nks05CRskC#DE0'H,oER#sCk'D0D2FI;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRRR--#kN0sCN0RoMCNP0HCR
RRRRRRRRRRRRRskC#D:0R=FRM0NR#0Nks05CRskC#DE0'H,oER#sCk'D0D2FI;R
RRRRRRRRRRMRC8VRH;R
RRRRRRRRRR-R-R#CDCCRs0MksR5jRHkMb0NRI#2Rj
RRRRRRRRCRRMH8RVR;
RRRRRRRRRR--CCD#R0sCkRsMjIR5s2Nb
RRRRRRRR8CMR;HV
RRRRCRRDV#HRs5NooEHERR>D0CV_8HMCRG20MEC
RRRRRRRRRHV5PHMCNO5sHoEoRE2=jR''02RE
CMRRRRRRRRRCRs8CkO8=R:RRFs5_0F#PkD5PHMCNO5sHoEo4E-RI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8C2;22
RRRRRRRRHRRVPRFCDsVF#I_0C$DRV=RH8GC_0#Nk0sNCMRN8CRs8CkO8RR='R4'0MEC
RRRRRRRRRRRRR--#kN0sCN0R#bFHP0HCR
RRRRRRRRRRCRs#0kDRR:=#kN0sCN0RC5s#0kD'oEHEs,RCD#k0F'DI
2;RRRRRRRRRDRC#RC
RRRRRRRRRHRRVsR5H0oE_8HMC>GRRoNsD2FIRC0EMR
RRRRRRRRRRRRRskC#DR0RRRRRR:RR=MRHPRCO5VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRRRRRRRRRMRRC#C8_ksFMM8Ho=R:RF5sk_M8#D0$CRR=VCHG8F_sk2M8;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRR#sCkRD05VDC0M_H8RCG8MFI0NFRsFoDI:2R=R
RRRRRRRRRRRRRRMRHPRCO5VDC0M_H8RCG8MFI0NFRsFoDI
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRR8sCk8OCRR:=NRM85_0F#PkD5PHMCNO5sHoEo4E-RI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8G222;R
RRRRRRRRRHFVRPVCsD_FI#D0$CRR=VCHG8N_#0Nks0NCRMs8RCO8kC=8RR''jRC0EMR
RRRRRRRRRRCRs#0kDRR:=MRF0#kN0sCN0RC5s#0kD'oEHEs,RCD#k0F'DI
2;RRRRRRRRRDRC#RC
RRRRRRRRRHRRVsR5H0oE_8HMC>GRRoNsD2FIRC0EMR
RRRRRRRRRRRRRskC#DR0RRRRRR:RR=MRHPRCO5VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2
RRRRRRRRRRRRMRRC#C8_ksFMM8Ho=R:RF5sk_M8#D0$CRR=VCHG8F_sk2M8;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRR#sCkRD05VDC0M_H8RCG8MFI0NFRsFoDI:2R=R
RRRRRRRRRRRRRRMRHPRCO5VDC0M_H8RCG8MFI0NFRsFoDI
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R
RRRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RoNsEEHoRR<=HCM0oRCsI0H8ER
RRRRRRVRHRs5NoIDFRR>=sEHo0M_H82CGRC0EMR
RRRRRRRRRskC#D50RNEsoHRoE8MFI0NFRsFoDI:2R=MRHP;CO
RRRRRRRR#CDCR
RRRRRRRRRskC#D50RNEsoHRoE8MFI0sFRH0oE_8HMCRG2:R=
RRRRRRRRRHRRMOPCRs5NooEHEFR8IFM0RosHEH0_MG8C2R;
RRRRRRRRRCMC8s#_F8kMHRMo:5=RsMFk80_#$RDC=HRVG_C8sMFk8R2;RR--sMFk8R
RRRRRRMRC8VRH;R
RRRRRRVRHRC5DVH0_MG8CRN>RsHoEoRE20MECR-R-Ro#HMGRC08CM
RRRRRRRRsRRCD#k0C5DVH0_MG8CRI8FMR0FNEsoH+oE4:2R=FR50sEC#>R=RPHMCNO5sHoEo2E2;R
RRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRR-R-Rk)FMs8RCD#k0R
RRRRRH5VRM8CC#F_skHM8MRo20MEC
RRRRRRRR#sCkRD0:s=RF8kM_GVHC58RNRsoRRRRRRRRR=RR>CRs#0kD,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRlsCN8HMCRsRRRRR=H>RMOPCRH5so_E0HCM8G
-4RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0NFRsFoDI
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRRPVCsD_FI#D0$C>R=RCFPsFVDI0_#$2DC;R
RRRRRCRM8H
V;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFMsHC#x
C;
-RR-HR#xsC_CV#Rk0MOH#FM
-RR-ERaCR#CVOkM0MHF#FROl0bkCER0CHR#xVCRsRFlNNRb#8#CRsPNHDNLCNRMlRC8"x#HCC_s#R"
RR--aRECF$MDRsbN0VRFRH0E#NRPsLHNDkCR#RC8HH0R0R'##CHx,0RHRRH#MCCPsNRb#8#C
-RR-FR0RDNRFsICRPDCCsDRFHk0M
C3RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRR:aR17p_zmBtQ_Be a;m)RRRRR-RR-ER#HCV08CRPOs0F
RRRRx#HCC_s#RR:z h)1emp k7_VCHG8R2RRRRRRR--VRFs#CHxRDFM$R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMRRVIRRRR:hRQa  t)=R:RMlHC#R5H_xCs'C#D,FIRx#HCC_s#F'DIR2;RR--OON0EHRD0NCsDR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58R#CHx_#sC'VDC0FR8IFM0R2VI;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<RR4FNsRsDo'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRD
#CRRRRRCRs#0kDRR:=0kF_VCHG8NR5sRoRRRRRR=RR>sRNoR,
RRRRRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CR>R=Rx#HCC_s#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMC=GR>HR#xsC_CD#'F;I2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FkGVHC
8;
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRsoRRRRR1:Raz7_pQmtB _eB)am;RRRRRRR-#-RE0HVCP8RCFO0sR
RRHR#xsC_C:#RR)zh p1me_ 7#GVHCR82RRRRR-R-RsVFRx#HCMRFDR$
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRMOF#M0N0IRVRRRRRQ:Rhta  :)R=HRlM5CR#CHx_#sC'IDF,HR#xsC_CD#'F;I2R-R-R0ONODERHs0CN
D#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85x#HCC_s#C'DV80RF0IMFIRV2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<RRRFsN'soDoCM0<ERRR420MEC
RRRRsRRCs0kMqRh1
w;RRRRCCD#
RRRRsRRCD#k0=R:R_0F#GVHC58RNRsoRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8G=RR>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCG=#>RH_xCs'C#D2FI;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_H#VG;C8
R
RVOkM0MHFR_0FkGVHC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRh:Rq)azqRp;RRRRRRRRR-RR-MRH0CCosR
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-V-RF#sRHRxCF$MD
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0D
C2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRFROMN#0MV0RIRRRRRR:Q hatR ):l=RHRMC5x#HCC_s#F'DI#,RH_xCs'C#D2FI;-RR-NRO0ROEDCH0s#ND
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRH5#xsC_CD#'CRV08MFI0VFRI
2;RCRLo
HMRRRRH5VRskC#DD0'C0MoERR<402RE
CMRRRRRCRs0MksRzhqwR;
RCRRD
#CRRRRRCRs#0kDRR:=0kF_VCHG8NR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=#>RH_xCs'C#EEHo,R
RRRRRRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CRRRR=#>RH_xCs'C#D,FI
RRRRRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FkGVHC
8;
VRRk0MOHRFM0#F_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRQa  t)R;RRRRRRRRRR-R-R0HMCsoC
RRRRx#HCC_s#RRRRRRRRRRRRRRRRz:Rh1) m pe7V_#H8GC;-RR-FRVsHR#xFCRM
D$RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRMOF#M0N0IRVRRRRRQ:Rhta  :)R=HRlM5CR#CHx_#sC'IDF,HR#xsC_CD#'F;I2R-R-R0ONODERHs0CN
D#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85x#HCC_s#C'DV80RF0IMFIRV2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwq1;R
RRDRC#RC
RRRRR#sCkRD0:0=RFV_#H8GCRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>HR#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_VCHG8
;
RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRq) pR;RR-RR-CRsNRD
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;RR--VRFs#CHxRDFM$R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02-RR-RRyFoVRk8NsR0LH#R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRO#FM00NMRRVIRRRR:hRQa  t)=R:RMlHC#R5H_xCs'C#D,FIRx#HCC_s#F'DIR2;RR--OON0EHRD0NCsDR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58R#CHx_#sC'VDC0FR8IFM0R2VI;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;zw
RRRR#CDCR
RRRRRskC#D:0R=FR0_HkVGRC85oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=Rx#HCC_s#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=Rx#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRRRRRkRoN_s8L#H0RRRRRR=>oskN8H_L0
#,RRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0kF_VCHG8
;
RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRq) pR;RR-RR-CRsNRD
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--VRFs#CHxRDFM$R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DC
RRRRMOF#M0N0kRoN_s8L#H0RRRRRh:Rq)azqRpRRRRRRRRRRRRRRRRRRR:=VCHG8k_oN_s8L#H02-RR-RRyFoVRk8NsR0LH#R
RRCRs0MksR)zh p1me_ 7#GVHCR8
R
H#RRRRO#FM00NMRRVIRRRR:hRQa  t)=R:RMlHC#R5H_xCs'C#D,FIRx#HCC_s#F'DIR2;RR--OON0EHRD0NCsDR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58R#CHx_#sC'VDC0FR8IFM0R2VI;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0shMRq;1w
RRRR#CDCR
RRRRRskC#D:0R=FR0_H#VGRC85oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRDRRC_V0HCM8GRRRR>R=Rx#HCC_s#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=Rx#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRRRRRkRoN_s8L#H0RRRRRR=>oskN8H_L0
#,RRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_VCHG8
;
RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;-RR-MRk#MHoCR8
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;R-RR-FRVsHR#xFCRM
D$RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRMOF#M0N0IRVRRRRRQ:Rhta  :)R=HRlM5CR#CHx_#sC'IDF,HR#xsC_CD#'F;I2R-R-R0ONODERHs0CN
D#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85x#HCC_s#C'DV80RF0IMFIRV2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<RRRFsN'soDoCM0<ERRR420MEC
RRRRsRRCs0kMqRhz
w;RRRRCCD#
RRRRsRRCD#k0=R:R_0FkGVHC58RNRsoRRRRRRRRR=RR>sRNoR,
RRRRRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>#CHx_#sC'IDF,R
RRRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRFRRPVCsD_FI#D0$C>R=RCFPsFVDI0_#$2DC;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_HkVG;C8

RRRkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 71hQt R7;RR--#MHoCR8
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHCR8;RR--VRFs#CHxRDFM$R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$2DC
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0VRIRR:RRRaQh )t RR:=lCHMRH5#xsC_CD#'FRI,#CHx_#sC'IDF2R;R-O-RNE0OR0DHCDsN#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8#R5H_xCs'C#D0CVRI8FMR0FV;I2
LRRCMoH
RRRRRHV5#sCk'D0DoCM0<ERRF4RssRNoC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwq1;R
RRDRC#RC
RRRRR#sCkRD0:0=RFV_#H8GCRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>HR#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$C
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_VCHG8
;
RkRVMHO0FsMRCx#HC
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-RbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;RR--VRFs#CHxRDFM$R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$2DC
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RORRF0M#NRM0VRIRR:RRRaQh )t RR:=lCHMRH5#xsC_CD#'FRI,#CHx_#sC'IDF2R;R-O-RNE0OR0DHCDsN#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp k7_VCHG8#R5H_xCs'C#EEHoRI8FMR0FV;I2
LRRCMoH
RRRRRHV5#sCk'D0DoCM0<ERRF4RssRNoC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhwqz;R
RRDRC#RC
RRRRR#sCkRD0:s=RCx#HCNR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRsRRH0oE_8HMCRGRR>R=Rx#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR#sCH;xC
R
RVOkM0MHFR#sCHRxC5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;R-H-RM0bk
RRRRx#HCC_s#RRRRRRRRRRRRRRRRz:Rh1) m pe7V_#H8GC;-RR-FRVsHR#xFCRM
D$RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DC
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRMOF#M0N0IRVRRRRRQ:Rhta  :)R=HRlM5CR#CHx_#sC'IDF,HR#xsC_CD#'F;I2R-R-R0ONODERHs0CN
D#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _H#VGRC85x#HCC_s#H'Eo8ERF0IMFIRV2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<RRRFsN'soDoCM0<ERRR420MEC
RRRRsRRCs0kMqRh1
w;RRRRCCD#
RRRRsRRCD#k0=R:R#sCHRxC5oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRosHEH0_MG8CRRRR=#>RH_xCs'C#D,FI
RRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D=CR>PRFCDsVF#I_0C$D2R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0FsMRCx#HC
;
R-R-RCmPsNDF8RC8lEN0RMVkOF0HMV#RFssRC
NDRkRVMHO0F"MR+5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MRDRR+0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs+R2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MRDRR+0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs+R2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR-5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MRDRR-0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM-R""
;
RkRVMHO0F"MR-5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs-R2R;
R8CMRMVkOF0HM-R""
;
RkRVMHO0F"MR-5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MRDRR-0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM-R""
;
RkRVMHO0F"MR-5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs-R2R;
R8CMRMVkOF0HM-R""
;
RkRVMHO0F"MR*5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MRDRR*0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM*R""
;
RkRVMHO0F"MR*5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs*R2R;
R8CMRMVkOF0HM*R""
;
RkRVMHO0F"MR*5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MRDRR*0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM*R""
;
RkRVMHO0F"MR*5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs*R2R;
R8CMRMVkOF0HM*R""
;
RkRVMHO0F"MR/5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MRDRR/0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MR/5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs/R2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MR/5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs: R)q
p2RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MRDRR/0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MR/5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs/R2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MRs"ClRR5
RDRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRR5DsRCl0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HMsR"C;l"
R
RVOkM0MHFRC"sl5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRlsCR;s2
CRRMV8Rk0MOHRFM"lsC"
;
RkRVMHO0F"MRs"ClRR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRR5DsRCl0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HMsR"C;l"
R
RVOkM0MHFRC"sl5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRlsCR;s2
CRRMV8Rk0MOHRFM"lsC"
;
RkRVMHO0F"MRl"F8RR5
RDRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRR5DlRF80kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HMlR"F;8"
R
RVOkM0MHFRF"l85"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIR8lFR;s2
CRRMV8Rk0MOHRFM"8lF"
;
RkRVMHO0F"MRl"F8RR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRR5DlRF80#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HMlR"F;8"
R
RVOkM0MHFRF"l85"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIR8lFR;s2
CRRMV8Rk0MOHRFM"8lF"
;
R-R-RCmPsNDF8RC8lEN0RMVkOF0HMV#RFHsRMo0CC
s#RkRVMHO0F"MR+5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMDR5R0+RFV_kH8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFR""+;R

RMVkOF0HM+R""
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,j+2RR;s2
CRRMV8Rk0MOHRFM";+"
R
RVOkM0MHFR""+RR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5+DRR_0F#GVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MR+
";
VRRk0MOHRFM"R+"5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,2RjRs+R2R;
R8CMRMVkOF0HM+R""
;
R-R-RCmPsNDF8RC8VOkM0MHF#R
RVOkM0MHFR""-RR5
RDRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:hzqa)2qp
RRRR0sCkRsMz h)1emp k7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5-DRR_0FkGVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MR-
";
VRRk0MOHRFM"R-"5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,2RjRs-R2R;
R8CMRMVkOF0HM-R""
;
RkRVMHO0F"MR-5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMDR5R0-RFV_#H8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFR""-;R

RMVkOF0HM-R""
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,j-2RR;s2
CRRMV8Rk0MOHRFM";-"
R
R-m-RPDCsFCN88kRVMHO0F
M#RkRVMHO0F"MR*5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMDR5R0*RFV_kH8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFR""*;R

RMVkOF0HM*R""
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,j*2RR;s2
CRRMV8Rk0MOHRFM";*"
R
RVOkM0MHFR""*RR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5*DRR_0F#GVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MR*
";
VRRk0MOHRFM"R*"5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,2RjRs*R2R;
R8CMRMVkOF0HM*R""
;
R-R-RCmPsNDF8RC8VOkM0MHF#R
RVOkM0MHFR""/RR5
RDRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:hzqa)2qp
RRRR0sCkRsMz h)1emp k7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5/DRR_0FkGVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MR/
";
VRRk0MOHRFM"R/"5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,2RjRs/R2R;
R8CMRMVkOF0HM/R""
;
RkRVMHO0F"MR/5"R
RRRR:DRR)zh p1me_ 7#GVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMDR5R0/RFV_#H8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFR""/;R

RMVkOF0HM/R""
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,j/2RR;s2
CRRMV8Rk0MOHRFM";/"
R
RVOkM0MHFRC"sl5"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMDR5RlsCR_0FkGVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MRs"Cl;R

RMVkOF0HMsR"CRl"5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,2RjRlsCR;s2
CRRMV8Rk0MOHRFM"lsC"
;
RkRVMHO0F"MRs"ClRR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5sDRC0lRFV_#H8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFRC"sl
";
VRRk0MOHRFM"lsC"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,js2RCslR2R;
R8CMRMVkOF0HMsR"C;l"
R
RVOkM0MHFRF"l85"R
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMDR5R8lFR_0FkGVHC58RsD,R'oEHEj,R2
2;RMRC8kRVMHO0F"MRl"F8;R

RMVkOF0HMlR"FR8"5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,2RjR8lFR;s2
CRRMV8Rk0MOHRFM"8lF"
;
RkRVMHO0F"MRl"F8RR5
RDRRRz:Rh1) m pe7V_#H8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8#RH
LRRCMoH
RRRR0sCkRsM5lDRF08RFV_#H8GCR,5sRED'H,oER2j2;R
RCRM8VOkM0MHFRF"l8
";
VRRk0MOHRFM"8lF"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,jl2RFs8R2R;
R8CMRMVkOF0HMlR"F;8"
R
R-F-RPDCsFCN88VRkH8GCRlOFbCNsRMVkOF0HMI#RHR0EHCM0o
CsRkRVMHO0F"MR=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:hzqa)2qpRRRRRRRRRRRRRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0=RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR""=;R

RMVkOF0HM/R"=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:hzqa)2qpRRRRRRRRRRRRRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5RR/=0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM/R"=
";
VRRk0MOHRFM"">=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs:qRhaqz)pR2RRRRRRRRRRRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5>DR=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:hzqa)2qpRRRRRRRRRRRRRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5RR<=0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM<R"=
";
VRRk0MOHRFM"R>"5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRahqzp)q2RRRRRRRRRRRRRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MRDRR>0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM>R""
;
RkRVMHO0F"MR<5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:hzqa)2qpRRRRRRRRRRRRRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0<RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR""<;R

RMVkOF0HM?R"=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:hzqa)2qpRRRRRRRRRRRRRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?0=RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR="?"
;
RkRVMHO0F"MR?"/=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs:qRhaqz)pR2RRRRRRRRRRRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD/R?=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"=?/"
;
RkRVMHO0F"MR?">=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs:qRhaqz)pR2RRRRRRRRRRRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD>R?=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"=?>"
;
RkRVMHO0F"MR?"<=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs:qRhaqz)pR2RRRRRRRRRRRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD<R?=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"=?<"
;
RkRVMHO0F"MR?R>"5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRahqzp)q2RRRRRRRRRRRRRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5RR?>0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R">
";
VRRk0MOHRFM""?<RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs:qRhaqz)pR2RRRRRRRRRRRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD<R?R_0FkGVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?;<"
R
RVOkM0MHFRGlNHllkRR5
RDRRRz:Rh1) m pe7V_kH8GC;RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRsRR:hzqa)2qp
RRRR0sCkRsMz h)1emp k7_VCHG8#RH
LRRCMoH
RRRR0sCkRsMlHNGlRkl5RD,0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HMNRlGkHll
;
RkRVMHO0FlMRHlMHk5lR
RRRR:DRR)zh p1me_ 7kGVHCR8;RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRRRs:qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMHRlMkHllDR5,FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFMlHHMl;kl
R
R-h-Rq)azq0pRFVRkH8GC
VRRk0MOHRFM"R="5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI=2RR;s2
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRR/=s
2;RMRC8kRVMHO0F"MR/;="
R
RVOkM0MHFR=">"
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRR>=s
2;RMRC8kRVMHO0F"MR>;="
R
RVOkM0MHFR="<"
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRR<=s
2;RMRC8kRVMHO0F"MR<;="
R
RVOkM0MHFR"">RR5
RDRRRh:Rq)azq
p;RRRRsRR:z h)1emp k7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kM0R5FV_kH8GCR,5DREs'H,oERDs'FRI2>2Rs;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs<R2R;
R8CMRMVkOF0HM<R""
;
RkRVMHO0F"MR?R="5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2=R?R;s2
CRRMV8Rk0MOHRFM""?=;R

RMVkOF0HM?R"/R="5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2/R?=2Rs;R
RCRM8VOkM0MHFR/"?=
";
VRRk0MOHRFM"=?>"
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_kH8GCR,5DREs'H,oERDs'FRI2?R>=s
2;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<R="5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2<R?=2Rs;R
RCRM8VOkM0MHFR<"?=
";
VRRk0MOHRFM""?>RR5
RDRRRh:Rq)azq
p;RRRRsRR:z h)1emp k7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI?2R>2Rs;R
RCRM8VOkM0MHFR>"?"
;
RkRVMHO0F"MR?R<"5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2<R?R;s2
CRRMV8Rk0MOHRFM""?<;R

RMVkOF0HMNRlGkHll
R5RRRRDRR:hzqa);qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRGlNHllkRF50_HkVGRC85RD,sH'EoRE,sF'DIR2,s
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5R
RRRRD:qRhaqz)pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0szMRh1) m pe7V_kH8GCR
H#RCRLo
HMRRRRskC0slMRHlMHk5lR0kF_VCHG8DR5,'RsEEHo,'RsD2FI,2Rs;R
RCRM8VOkM0MHFRMlHHllk;R

RR--FsPCD8FNCk8RVCHG8FROlsbNCkRVMHO0FRM#IEH0RNsCDR
RVOkM0MHFR""=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs: R)q
p2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"
R5RRRRDRR:z h)1emp k7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5RR/=0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM/R"=
";
VRRk0MOHRFM"">=RR5
RDRRRz:Rh1) m pe7V_kH8GC;R
RRRRs: R)q
p2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D>0=RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR=">"
;
RkRVMHO0F"MR<R="5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRq) pR2
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5<DR=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM""<=;R

RMVkOF0HM>R""
R5RRRRDRR:z h)1emp k7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0>RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""
R5RRRRDRR:z h)1emp k7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0<RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR""<;R

RMVkOF0HM?R"=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:)p q2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5RR?=0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R"=
";
VRRk0MOHRFM"=?/"
R5RRRRDRR:z h)1emp k7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?R/=0kF_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R"/;="
R
RVOkM0MHFR>"?=5"R
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:)p q2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5R=?>R_0FkGVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<R="5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRq) pR2
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD<R?=FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"=?<"
;
RkRVMHO0F"MR?R>"5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRq) pR2
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD>R?R_0FkGVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?;>"
R
RVOkM0MHFR<"?"
R5RRRRDRR:z h)1emp k7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?0<RFV_kH8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR<"?"
;
RkRVMHO0FlMRNlGHk5lR
RRRR:DRR)zh p1me_ 7kGVHC
8;RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRGlNHllkR,5DR_0FkGVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5R
RRRRD:hRz)m 1p7e _HkVG;C8
RRRR:sRRq) pR2
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMHRlMkHllDR5,FR0_HkVGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFMlHHMl;kl
R
R-s-RCRNDNRM8kGVHCR8
RMVkOF0HM=R""
R5RRRRDRR:)p q;R
RRRRs:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2RR=s
2;RMRC8kRVMHO0F"MR=
";
VRRk0MOHRFM""/=RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRR/=s
2;RMRC8kRVMHO0F"MR/;="
R
RVOkM0MHFR=">"
R5RRRRDRR:)p q;R
RRRRs:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2=R>R;s2
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI<2R=2Rs;R
RCRM8VOkM0MHFR="<"
;
RkRVMHO0F"MR>5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI>2RR;s2
CRRMV8Rk0MOHRFM";>"
R
RVOkM0MHFR""<RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0kF_VCHG8DR5,'RsEEHo,'RsD2FIRs<R2R;
R8CMRMVkOF0HM<R""
;
RkRVMHO0F"MR?R="5R
RRRRD: R)q
p;RRRRsRR:z h)1emp k7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI?2R=2Rs;R
RCRM8VOkM0MHFR="?"
;
RkRVMHO0F"MR?"/=RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_kH8GCR,5DREs'H,oERDs'FRI2?R/=s
2;RMRC8kRVMHO0F"MR?"/=;R

RMVkOF0HM?R">R="5R
RRRRD: R)q
p;RRRRsRR:z h)1emp k7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_HkVGRC85RD,sH'EoRE,sF'DI?2R>s=R2R;
R8CMRMVkOF0HM?R">;="
R
RVOkM0MHFR<"?=5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_kH8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0FkGVHC58RDs,R'oEHEs,R'IDF2<R?=2Rs;R
RCRM8VOkM0MHFR<"?=
";
VRRk0MOHRFM""?>RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_kH8GCR,5DREs'H,oERDs'FRI2?s>R2R;
R8CMRMVkOF0HM?R">
";
VRRk0MOHRFM""?<RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_kH8GCR,5DREs'H,oERDs'FRI2?s<R2R;
R8CMRMVkOF0HM?R"<
";RRR
RMVkOF0HMNRlGkHll
R5RRRRDRR:)p q;R
RRRRs:hRz)m 1p7e _HkVG2C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMhRz)m 1p7e _HkVGRC8HR#
RoLCHRM
RsRRCs0kMNRlGkHll0R5FV_kH8GCR,5DREs'H,oERDs'F,I2R;s2
CRRMV8Rk0MOHRFMlHNGl;kl
R
RVOkM0MHFRMlHHllkRR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7kGVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRMlHHllkRF50_HkVGRC85RD,sH'EoRE,sF'DIR2,s
2;RMRC8kRVMHO0FlMRHlMHk
l;
-RR-PRFCFsDN88CRH#VGRC8ObFlNRsCVOkM0MHF#HRI0HERMo0CCRs
RMVkOF0HM=R""
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRRQ:Rhta  
)2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D=FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRRQ:Rhta  
)2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D/0=RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR="/"
;
RkRVMHO0F"MR>R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MRD=R>R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR>;="
R
RVOkM0MHFR="<"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRRQ:Rhta  
)2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D<0=RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR="<"
;
RkRVMHO0F"MR>5"R
RRRR:DRR)zh p1me_ 7#GVHC
8;RRRRsRR:Q hat2 )
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0>RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRRQ:Rhta  
)2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D<FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM";<"
R
RVOkM0MHFR="?"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRRQ:Rhta  
)2RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5?DR=FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM""?=;R

RMVkOF0HM?R"/R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5R=?/R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?"/=;R

RMVkOF0HM?R">R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5R=?>R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5R=?<R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?"<=;R

RMVkOF0HM?R">5"R
RRRR:DRR)zh p1me_ 7#GVHC
8;RRRRsRR:Q hat2 )
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?0>RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR>"?"
;
RkRVMHO0F"MR?R<"5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5RR?<0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R"<
";
VRRk0MOHRFMlHNGlRkl5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRGlNHllkR,5DR_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRMlHHllkR,5DR_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0FlMRHlMHk
l;
-RR-MRH0CCosMRN8VR#H8GC
VRRk0MOHRFM"R="5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI=2RR;s2
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRR/=s
2;RMRC8kRVMHO0F"MR/;="
R
RVOkM0MHFR=">"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRR>=s
2;RMRC8kRVMHO0F"MR>;="
R
RVOkM0MHFR="<"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRR<=s
2;RMRC8kRVMHO0F"MR<;="
R
RVOkM0MHFR"">RR5
RDRRRQ:Rhta  
);RRRRsRR:z h)1emp #7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kM0R5FV_#H8GCR,5DREs'H,oERDs'FRI2>2Rs;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs<R2R;
R8CMRMVkOF0HM<R""
;
RkRVMHO0F"MR?R="5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2=R?R;s2
CRRMV8Rk0MOHRFM""?=;R

RMVkOF0HM?R"/R="5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2/R?=2Rs;R
RCRM8VOkM0MHFR/"?=
";
VRRk0MOHRFM"=?>"
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_#H8GCR,5DREs'H,oERDs'FRI2?R>=s
2;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<R="5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2<R?=2Rs;R
RCRM8VOkM0MHFR<"?=
";
VRRk0MOHRFM""?>RR5
RDRRRQ:Rhta  
);RRRRsRR:z h)1emp #7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI?2R>2Rs;R
RCRM8VOkM0MHFR>"?"
;
RkRVMHO0F"MR?R<"5R
RRRRD:hRQa  t)R;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2<R?R;s2
CRRMV8Rk0MOHRFM""?<;R

RMVkOF0HMNRlGkHll
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0slMRNlGHk5lR0#F_VCHG8DR5,'RsEEHo,'RsD2FI,2Rs;R
RCRM8VOkM0MHFRGlNHllk;R

RMVkOF0HMHRlMkHll
R5RRRRDRR:Q hat; )
RRRR:sRR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0slMRHlMHk5lR0#F_VCHG8DR5,'RsEEHo,'RsD2FI,2Rs;R
RCRM8VOkM0MHFRMlHHllk;R

RR--FsPCD8FNC#8RVCHG8FROlsbNCkRVMHO0FRM#IEH0RNsCDR
RVOkM0MHFR""=RR5
RDRRRz:Rh1) m pe7V_#H8GC;R
RRRRs: R)q
p2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D=FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5RR/=0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM/R"=
";
VRRk0MOHRFM"">=RR5
RDRRRz:Rh1) m pe7V_#H8GC;R
RRRRs: R)q
p2RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRR5D>0=RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR=">"
;
RkRVMHO0F"MR<R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRq) pR2
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5<DR=FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM""<=;R

RMVkOF0HM>R""
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0>RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMDR5R0<RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR""<;R

RMVkOF0HM?R"=5"R
RRRR:DRR)zh p1me_ 7#GVHC
8;RRRRsRR:)p q2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5RR?=0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R"=
";
VRRk0MOHRFM"=?/"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?R/=0#F_VCHG8sR5,'RDEEHo,'RDD2FI2R;
R8CMRMVkOF0HM?R"/;="
R
RVOkM0MHFR>"?=5"R
RRRR:DRR)zh p1me_ 7#GVHC
8;RRRRsRR:)p q2R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMDR5R=?>R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<R="5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRq) pR2
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD<R?=FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFM"=?<"
;
RkRVMHO0F"MR?R>"5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRq) pR2
RsRRCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0s5MRD>R?R_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0F"MR?;>"
R
RVOkM0MHFR<"?"
R5RRRRDRR:z h)1emp #7_VCHG8R;
RsRRR):R 2qp
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRR5D?0<RFV_#H8GCR,5sRED'H,oERDD'F2I2;R
RCRM8VOkM0MHFR<"?"
;
RkRVMHO0FlMRNlGHk5lR
RRRR:DRR)zh p1me_ 7#GVHC
8;RRRRsRR:)p q2R
RRCRs0MksR)zh p1me_ 7#GVHCH8R#R
RLHCoMR
RRCRs0MksRGlNHllkR,5DR_0F#GVHC58RsD,R'oEHED,R'IDF2
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5R
RRRRD:hRz)m 1p7e _H#VG;C8
RRRR:sRRq) pR2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMHRlMkHllDR5,FR0_H#VGRC85Rs,DH'EoRE,DF'DI;22
CRRMV8Rk0MOHRFMlHHMl;kl
R
R-)-R RqpNRM8#GVHCR8
RMVkOF0HM=R""
R5RRRRDRR:)p q;R
RRRRs:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2RR=s
2;RMRC8kRVMHO0F"MR=
";
VRRk0MOHRFM""/=RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRR/=s
2;RMRC8kRVMHO0F"MR/;="
R
RVOkM0MHFR=">"
R5RRRRDRR:)p q;R
RRRRs:hRz)m 1p7e _H#VG2C8RRRRRRRRRRRRR-R-RGVHCb8RF0HMRbHMkR0
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2=R>R;s2
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI<2R=2Rs;R
RCRM8VOkM0MHFR="<"
;
RkRVMHO0F"MR>5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI>2RR;s2
CRRMV8Rk0MOHRFM";>"
R
RVOkM0MHFR""<RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s5MR0#F_VCHG8DR5,'RsEEHo,'RsD2FIRs<R2R;
R8CMRMVkOF0HM<R""
;
RkRVMHO0F"MR?R="5R
RRRRD: R)q
p;RRRRsRR:z h)1emp #7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI?2R=2Rs;R
RCRM8VOkM0MHFR="?"
;
RkRVMHO0F"MR?"/=RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_#H8GCR,5DREs'H,oERDs'FRI2?R/=s
2;RMRC8kRVMHO0F"MR?"/=;R

RMVkOF0HM?R">R="5R
RRRRD: R)q
p;RRRRsRR:z h)1emp #7_VCHG8R2RRRRRRRRRRRRR-V-RH8GCRHbFMH0RM0bk
RRRR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRF50_H#VGRC85RD,sH'EoRE,sF'DI?2R>s=R2R;
R8CMRMVkOF0HM?R">;="
R
RVOkM0MHFR<"?=5"R
RRRR:DRRq) pR;
RsRRRz:Rh1) m pe7V_#H8GC2RRRRRRRRRRRR-RR-HRVGRC8bMFH0MRHb
k0RRRRskC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsM5_0F#GVHC58RDs,R'oEHEs,R'IDF2<R?=2Rs;R
RCRM8VOkM0MHFR<"?=
";
VRRk0MOHRFM""?>RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_#H8GCR,5DREs'H,oERDs'FRI2?s>R2R;
R8CMRMVkOF0HM?R">
";
VRRk0MOHRFM""?<RR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHCR82RRRRRRRRRRRRRR--VCHG8FRbHRM0HkMb0R
RRCRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kM0R5FV_#H8GCR,5DREs'H,oERDs'FRI2?s<R2R;
R8CMRMVkOF0HM?R"<
";
VRRk0MOHRFMlHNGlRkl5R
RRRRD: R)q
p;RRRRsRR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMNRlGkHll0R5FV_#H8GCR,5DREs'H,oERDs'F,I2R;s2
CRRMV8Rk0MOHRFMlHNGl;kl
R
RVOkM0MHFRMlHHllkRR5
RDRRR):R ;qp
RRRR:sRR)zh p1me_ 7#GVHC
82RRRRskC0szMRh1) m pe7V_#H8GCR
H#RCRLo
HMRRRRskC0slMRHlMHk5lR0#F_VCHG8DR5,'RsEEHo,'RsD2FI,2Rs;R
RCRM8VOkM0MHFRMlHHllk;-

-sRbNNolRM#$0#ECHF#_V-V
-0RsD$_#MC0E#RH#F
VV
-RR-FROb8HCRFVsl0R#8F_Do_HO00CGHRF
Rb0$CeRvpDgbkH#R#'R5zR',',X'R''j,4R''',RZR',',W'R''p,]R''',R-R',CFsss
2;R$R0bOCRE_NsHCM8G_C8Lv$_eRpgHN#Rs$sNRa517p_zmBtQ2VRFRqB])aqB 
);R$R0bvCRe_pgHCM8G_C8LO$_ERNsHN#Rs$sNR]5BqB)qa2 )RRFV1_a7ztpmQ
B;R$R0bvCRebpgD_k#HCM8G_C8LO$_ERNsHN#Rs$sNR]5BqB)qa2 )RRFVvgepb#Dk;R

RMOF#M0N0eRvp0g_FE_ON:sRRNOEsM_H8CCG8$_L_pveg=R:RX"zjW4Zp"]-;R
RO#FM00NMRNOEsF_0_pvegRR:vgep_8HMC8GC__L$OsENR
:=RRRR5''zRR=>',z'R''XRR=>',X'R''jRR=>',j'R''4RR=>',4'R''ZRR=>',Z'
RRRRWR''>R=R''W,pR''>R=R''p,]R''>R=R''],-R''>R=R''-,0RFE#CsRR=>'2z';R
RO#FM00NMRNOEsF_0_pvegkbD#RR:vgepb#Dk_8HMC8GC__L$OsENR
:=RRRR5''zRR=>',z'R''XRR=>',X'R''jRR=>',j'R''4RR=>',4'R''ZRR=>',Z'
RRRRWR''>R=R''W,pR''>R=R''p,]R''>R=R''],-R''>R=R''-,0RFE#CsRR=>CFsss
2;RFROMN#0Mh0RAR1u:]RBqB)qaR )RRRRRR:=B)]qq Ba)N'PDn54jR2;RR--#ObNCERONOsN0
CsRFROMN#0Mh0RzR1R:aR1)tQh50.RF2R4RR:=5EF0CRs#='>RR;'2

RRR-R-RsbkbCF#:	R1HRb#I0EHCbR#N
OCRsRbF8OCkRsC#b	H_HIE0bC#NROC5R
RRRRp:MRHFRk0p Qh2#RH
RRRRsPNHDNLCCRsN	8mRA:Rm mpq
h;RRRRPHNsNCLDR:ORRqB])aqB 
);RCRLo
HMRRRRIDEHCRRp/M=RkRDDNRM8pD3NDC'DMEo0RR/=jFRDFRb
RRRRRRHV5Np3D4D52RR='RR'FpsR3DND5R42=ARh1FuRs3RpN5DD4=2RR2]aRC0EMR
RRRRRRCRsN58RDO,R,CRsN	8m2R;
RRRRR#CDCR
RRRRRRGRCH
0;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RMRC8sRbF8OCkRsC#b	H_HIE0bC#N;OC
R
R-b-RkFsb#RC:I0sHCV#RH8GCRHbFMH0RMR0FNHRDMRC
RFbsOkC8sICRsCH0RR5
RpRRRRRRRRRRRH:RM0FkRhpQ R;RRRRRRRRRRRRRRR--HkMb0HRDMRC
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7kGVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RH
RRRRsPNHDNLCRR#RRRR:aR1)tQh504RFNRPD'kCDoCM0+ER4:2R=FR50sEC#>R=R''R2R;
RPRRNNsHLRDC#8HMGRR:Q hat; )
LRRCMoHR-R-RMVkOF0HMsRIHR0CRGR NDlbCj:Rj3444j4j
RRRRM#H8:GR=;R4
RRRRsVFRHHRMNRPD'kCEEHoRI8FMR0FPkNDCF'DIFRDFRb
RRRRRRHVHRR=-04RE
CMRRRRRRRR#H5#M28GRR:=';3'
RRRRRRRRM#H8RGRR=R:RM#H8+GRR
4;RRRRRMRC8VRH;R
RRRRR#H5#M28GRR:=vgep__0FOsEN571a_mzpt5QBPkNDC25H2
2;RRRRRHR#MR8GR:RR=HR#MR8G+;R4
RRRR8CMRFDFbR;
RIRRsCH05RD,#[,RkH#0V8HC,HRVC2D8;R
RCRM8bOsFCs8kCsRIH;0C
R
R-b-RkFsb#RC:I0sHCV#RH8GCRHbFMH0RMR0FNHRDMRC
RFbsOkC8sICRsCH0RR5
RpRRRRRRRRRRRH:RM0FkRhpQ R;RRRRRRRRRRRRRRR--HkMb0HRDMRC
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7#GVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RH
RRRRsPNHDNLCRR#RRRR:aR1)tQh504RFNRPD'kCDoCM0+ER4
2;RRRRPHNsNCLDRM#H8:GRRaQh )t ;R
RLHCoM-RR-kRVMHO0FIMRsCH0R RRGbNlDRC:j4j43j44jR
RRHR#MR8G:4=R;R
RRFRVsRRHHPMRNCDk'oEHEFR8IFM0RDPNkDC'FDIRF
FbRRRRRVRHR=HRRR-40MEC
RRRRRRRR##5HGM82=R:R''3;R
RRRRRRHR#MR8GR:RR=HR#MR8G+;R4
RRRRCRRMH8RVR;
RRRRR##5HGM82=R:RpvegF_0_NOEsa517p_zmBtQ5DPNkHC52;22
RRRR#RRHGM8RRRR:#=RHGM8R4+R;R
RRMRC8FRDF
b;RRRRI0sHC,5DRR#,[0k#HCVH8V,RH8CD2R;
R8CMRFbsOkC8sICRsCH0;R

RFbsOkC8s)CR 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_kH8GC2#RH
RRRRR--u#F#HCLDR08NNR:Rjjjjjj3jjjjjjR
RR-R-RRRRRRRRRRRRRRRRRjjjjjjjjjjjjR
RRNRPsLHNDOCRRRRRRRR:B)]qq Ba)R;
RPRRNNsHLRDCs8CNm:	RRmAmph q;R
RRNRPsLHNDHCRRRRRRRR:Q hat; )RRRRRRRRR-R-R8HMCPGRNNsHL
DCRRRRPHNsNCLDRRlP:VRkH8GCRq5ep'z soNMC
2;RRRRPHNsNCLDR#DN0RkR:mRAmqp h=R:RDVN#RC;RRRRR-R-R#DN0ERONOsN0RCsIRN#N"MR_R"
RPRRNNsHLRDCVMFk808FRA:Rm mpq:hR=NRVD;#CR-R-RkVFMN8RR""3
LRRCMoHR-R-Rq) 7R
RRqRepRz :5=Rezqp N'sMRoC='>Rz;'2
RRRRH1	bE_IH#0CbCNOR25p;R
RRVRHRpeqzD 'C0MoERR>jER0CRMRRRRRRRRRR-R-RMMFRDhkDMRHbRk0#H0sMRo
RRRRRNsC8DR5,,RORNsC82m	;R
RRRRRH=R:RDPNkEC'H;oE
RRRRIRRECHDR>HR=qRep'z DRFIDbFF
RRRRRRRRRHVs8CNm=	RRDVN#0CRERCMRRRRRRRRRRRRRR--ADNHR0FkRRHV0sECCNRI#RRNLRN8s8CN
RRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCRR&"q) 7V5kH8GC2
R"RRRRRRRRRRRR& R"MF8RV0R#soHMROCMF0kMC8sC"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s
M;RRRRRRRRCHD#VRRO=_R''ER0CRM
RRRRRRRRRRHVHRR=PkNDCH'Eo0ERE
CMRRRRRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_Ml&CRR ")qk75VCHG8"2R
RRRRRRRRRRRR&RRR0"1soHMRoLCHRM#IEH0RRNM"""_"#"RCsPCHR0$CFsssR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR#CDHDVRNk#0RC0EMR
RRRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNlR"&R)7 q5HkVG2C8RR"
RRRRRRRRRRRRR"&RaRIFkCM8sF#OsRC#8CC0O80CRRHMHkMb00R#soHMR_""_"""
RRRRRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR#CDCR
RRRRRRRRRRNRD#R0k:0=Rs;kC
RRRRRRRRCRRMH8RVR;
RRRRRCRRDV#HR=ORR''3RC0EMRRRRRRRRRRRRRRRRR--LNHMsb$RF0HM
RRRRRRRRHRRVFRVk8M8F00RE
CMRRRRRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_Ml&CRR ")qk75VCHG8"2R
RRRRRRRRRRRR&RRRI"aFHRLM$NsRHbFMR0#VMFk8MRHRbHMk#0R0MsHo#"RCsPCHR0$CFsssR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR#CDHHVRRR/=-04RERCMRRRRRRRRRRRRRRRR-1-RCsbCNs0FRRHM0RECIMsFobR#FR0
RRRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCRR&"q) 7V5kH8GC2
R"RRRRRRRRRRRRRRR&"O7CHDlNRHbFM80RFRC#MRF0lON0EkRMlsLCRsVFlRN0"R
RRRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRRRRskC0s
M;RRRRRRRRRMRC8VRH;R
RRRRRRRRRVMFk808FRR:=0Csk;R
RRRRRRRRRD0N#k=R:RDVN#
C;RRRRRRRRCHD#VRRO=RR''sRFR=ORR1hAusRFR=ORRR]a0MECR-R-RNsC8oHMRM8FCR3
RRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_NRlC&)R" 5q7kGVHCR82"R
RRRRRRRRRRRR&"F1Ess0RC,N8RN1bOCCRMkOFM80CRRHMHkMb00R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s
M;RRRRRRRRCHD#VERON0s_Fe_vpDgbkO#52RR=CFsssER0CRM
RRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_NRlC&)R" 5q7kGVHCR82"R
RRRRRRRRRRRR&"NBEs0NOC'sR"
R&RRRRRRRRRRRRORR&"s'RC,N8RbCGCCO08aR17p_zmBtQR0DHCDsN3R"
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCk;sM
RRRRRRRR#CDCR
RRRRRRRRRlHP52=R:RNOEsF_0_pveg25O;R
RRRRRRRRRH=R:R-HRR
4;RRRRRRRRRVRHR<HRR'lPDRFI0MEC
RRRRRRRRRRRRpeqz: R=PRl;R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCRM8H
V;RRRRRRRRRNRD#R0k:V=RNCD#;R
RRRRRRMRC8VRH;R
RRRRRRCRsNp85,,RORNsC82m	;R
RRRRRCRM8DbFF;R
RRMRC8VRH;R
RCRM8bOsFCs8kC R)q
7;
bRRsCFO8CksRq) 7R5pRRRR:MRHFRk0p Qh;R
RRRRRRRRRRRRRReRRq pzRF:RkR0RR)zh p1me_ 7kGVHC
8;RRRRRRRRRRRRRRRRRmtm7:RRR0FkRARRm mpqRh2HR#
R-RR-FRu#L#HD8CRN:0NRjRjj3jjjjjjj
jjRRRR-R-RRRRRRRRRRRRRRjRRjjjjjjjjj
jjRRRRPHNsNCLDRRORRRRR:]RBqB)qa; )
RRRRsPNHDNLCCRsN	8mRA:Rm mpq
h;RRRRPHNsNCLDRRlP:VRkH8GCRq5ep'z soNMC
2;RRRRPHNsNCLDRRHRRRRR:hRQa  t)R;RRRRRRRRR-H-RMG8CRsPNHDNLCR
RRNRPsLHNDDCRNk#0RRR:Apmm Rqh:V=RNCD#;RRRRRRR-D-RNR#0OsENNCO0sNRI#MRNR""_
RRRRsPNHDNLCFRVk8M8F:0RRmAmph qRR:=V#NDCR;R-V-RF8kMR"NR3R"
RoLCHRMR-)-R 
q7RRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;
R1RR	_HbI0EHCN#bO5CRp
2;RRRRHeVRq pz'MDCoR0E>RRj0MEC
RRRRsRRCRN85RD,Os,RCmN8	
2;RRRRRRRH:P=RNCDk'oEHER;
RRRRRmtm7=R:RDVN#
C;RRRRRERIHRDCH=R>RpeqzD 'FDIRF
FbRRRRRRRRHMVRFs0RCmN8	ER0CRMRR-RR-NRAHFDRkH0RVER0CRsCIRN#NNRL8CRsNR8
RRRRRRRRR0sCk;sM
RRRRRRRR#CDHOVRR'=R_0'RE
CMRRRRRRRRRVRHR=HRRDPNkEC'HRoE0MECRRRRRRRRR-R-RoACHRM#IEH0RRNM"
_"RRRRRRRRRRRRskC0s
M;RRRRRRRRRDRC#RHVD0N#kER0CRMRRRRRRRRRRRRRRR--""__R08CCCO08R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCCD#
RRRRRRRRRRRR#DN0:kR=sR0k
C;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVORR='R3'0MECRRRRRRRRRRRRRRRR-L-RHsMN$FRbH
M0RRRRRRRRRVRHRkVFMF880ER0CRM
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR#CDHHVRRR/=-04RERCMRRRRRRRRRRRRRRRR-1-RCsbCNs0FRRHM0RECIMsFobR#FR0
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR8CMR;HV
RRRRRRRRVRRF8kM8RF0:0=Rs;kC
RRRRRRRRDRRNk#0RR:=V#NDCR;
RRRRRCRRDV#HRE5ON0s_Fe_vpDgbkO#52RR=CFsss02RERCMR-R-RDQDCDoNRNOEs0NOC#s/E0FsRNsC8R
RRRRRRRRRskC0s
M;RRRRRRRRCCD#
RRRRRRRRlRRP25HRR:=OsEN__0Fvgep5;O2
RRRRRRRRHRRRR:=HRR-4R;
RRRRRRRRRRHVHRR<lDP'F0IRERCMRRRRRRRRRRRR-s-RCHN8M8oRF
MCRRRRRRRRRRRRt7mmRR:=0Csk;R
RRRRRRRRRRqRepRz :l=RPR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR8CMR;HV
RRRRRRRRDRRNk#0RR:=V#NDCR;
RRRRRCRRMH8RVR;
RRRRRsRRC5N8pO,R,CRsN	8m2R;
RRRRR8CMRFDFbR;
RCRRD
#CRRRRRmRtm:7R=sR0kRC;RRRRRRRRRRRRRRRRR-R-RNsC8MRH0NFRRDMkDsRNs
N$RRRRCRM8H
V;RMRC8sRbF8OCkRsC)7 q;R

RFbsOkC8s)CR 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_#H8GC2#RH
RRRRsPNHDNLCRRORRRRRB:R]qq)B)a ;R
RRNRPsLHNDsCRCmN8	RR:Apmm ;qh
RRRRsPNHDNLCRRHRRRRRQ:Rhta  R);RRRRRRRRRR--HCM8GNRPsLHNDRC
RPRRNNsHLRDCl:PRRH#VGRC85peqzs 'NCMo2R;
RPRRNNsHLRDCD0N#k:RRRmAmph qRR:=V#NDCR;RRRRRRR--D0N#RNOEs0NOCIsRNN#RM_R""R
RRNRPsLHNDVCRF8kM8RF0:mRAmqp h=R:RDVN#RC;RR--VMFk8RRN"
3"RCRLoRHMRR--)7 q
RRRRpeqz: R=eR5q pz'MsNo=CR>zR''
2;RRRR1b	H_HIE0bC#NROC5;p2
RRRRRHVezqp C'DMEo0Rj>RRC0EMRRRRRRRRRRRRR--MRFMhDkDRbHMk#0R0MsHoR
RRRRRs8CNR,5DRRO,s8CNm;	2
RRRRHRRRR:=PkNDCH'Eo
E;RRRRRERIHRDCH=R>RpeqzD 'FDIRF
FbRRRRRRRRHsVRCmN8	RR=V#NDCER0CRMRRRRRRRRRRRRR-A-RNRHDFRk0H0VRECCsR#INRLNRNs8RC
N8RRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNlR"&R)7 q5H#VG2C8RR"
RRRRRRRRR&RRRM" 8VRFRs#0HRMoCFMOkCM0s"C8
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRDV#HR=ORR''_RC0EMR
RRRRRRRRRHHVRRP=RNCDk'oEHEER0CRM
RRRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCRR&"q) 7V5#H8GC2
R"RRRRRRRRRRRRRRR&"s10HRMoLHCoMI#RHR0EN"MR""_""CR#PHCs0C$RsssF;R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCHD#VNRD#R0k0MEC
RRRRRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_NRlC&)R" 5q7#GVHCR82"R
RRRRRRRRRRRRR&aR"IkFRMs8C#sOFC8#RCO0C0RC8HHMRM0bkRs#0HRMo"_"_"
""RRRRRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCCD#
RRRRRRRRRRRR#DN0:kR=sR0k
C;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVORR='R3'0MECRRRRRRRRRRRRRRRR-L-RHsMN$FRbH
M0RRRRRRRRRVRHRkVFMF880ER0CRM
RRRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCRR&"q) 7V5#H8GC2
R"RRRRRRRRRRRRRRR&"FaIRMLHNRs$bMFH0V#RF8kMRRHMHkMb00R#soHM"CR#PHCs0C$RsssF;R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCHD#VRRH/-=R4ER0CRMRRRRRRRRRRRRRR-RR-CR1bNCs0RFsH0MREICRsoFMRF#b0R
RRRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNlR"&R)7 q5H#VG2C8RR"
RRRRRRRRRRRRR"&R7HCOlRNDbMFH0FR8CM#RFl0RNE0ORlMkLRCsVlFsN"0R
RRRRRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR8CMR;HV
RRRRRRRRVRRF8kM8RF0:0=Rs;kC
RRRRRRRRDRRNk#0RR:=V#NDCR;
RRRRRCRRDV#HR=ORR''RRRFsORR=huA1RRFsORR=]0aRERCMRR--s8CNHRMo8CFM3R
RRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_Ml&CRR ")q#75VCHG8"2R
RRRRRRRRRRRR"&R1sEF0CRsNR8,1ObNCMRCOMFk0RC8HHMRM0bkRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRDV#HRNOEsF_0_pvegkbD#25ORC=RsssFRC0EMR
RRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_Ml&CRR ")q#75VCHG8"2R
RRRRRRRRRRRR"&RBsENNCO0s"R'RR&
RRRRRRRRRORRR"&R'CRsNR8,CCGbO80CR71a_mzptRQBDCH0s3ND"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s
M;RRRRRRRRCCD#
RRRRRRRRlRRP25HRR:=OsEN__0Fvgep5;O2
RRRRRRRRHRRRR:=HRR-4R;
RRRRRRRRRRHVHRR<lDP'F0IRE
CMRRRRRRRRRRRRezqp =R:R;lP
RRRRRRRRRRRR0sCk;sM
RRRRRRRRCRRMH8RVR;
RRRRRRRRR#DN0:kR=NRVD;#C
RRRRRRRR8CMR;HV
RRRRRRRRNsC8,5pRRO,s8CNm;	2
RRRRCRRMD8RF;Fb
RRRR8CMR;HV
CRRMb8RsCFO8CksRq) 7
;
RsRbF8OCkRsC)7 q5RpRR:RRRFHMkp0RQ;h 
RRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp #7_VCHG8R;
RRRRRRRRRRRRRRRRt7mmRRR:FRk0RmRAmqp hH2R#R
RRNRPsLHNDPCRNCDk_HkVGRC8:hRz)m 1p7e _HkVGRC85peqzs 'NCMo2R;
RoLCHRMR-)-R 
q7RRRR)7 qRR5p=p>R,qRepRz =P>RNCDk_HkVG,C8Rmtm7>R=Rmtm7
2;RRRRezqp =R:R)zh p1me_ 7#GVHC58RPkNDCV_kH8GC2R;
R8CMRFbsOkC8s)CR ;q7
R
R-F-ROD0NRNsC8MRN8sRIH
0CRsRbF8OCkRsCFHIs05CR
RRRRRpRRRRRR:RRRFHMkp0RQ;h RRRRRRRRRRRRR-RR-MRHbRk0DCHM
RRRRpeqzR RR:RRRRHMRzRRh1) m pe7V_kH8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRKaz1Q wQ7RR:HRMRRQR17R R:s=RH0oE;R
RRQRw Rp7RRRR:MRHRRRRWaQ7]=R:RRj2HR#
RoLCHRMR- -RGbNlDjCRdj3d
RRRRHIs05CRpRRRRRRRR>R=R
p,RRRRRRRRReRRq pzRRRRRR=>0FF_#H0sM5oRezqp 
2,RRRRRRRRRKRRzQ1aw7Q RR=>Kaz1Q wQ7R,
RRRRRRRRRQRw Rp7RRRR=w>RQ7 p2R;
R8CMRFbsOkC8sFCRI0sHC
;
RsRbF8OCkRsCFHIs05CR
RRRRRpRRRRRR:RRRFHMkp0RQ;h RRRRRRRRRRRRR-RR-MRHbRk0DCHM
RRRRpeqzR RR:RRRRHMRzRRh1) m pe7V_#H8GC;-RR-HRVGRC8bMFH0MRHb
k0RRRRKaz1Q wQ7RR:HRMRRQR17R R:s=RH0oE;R
RRQRw Rp7RRRR:MRHRRRRWaQ7]=R:RRj2HR#
RoLCHRMR- -RGbNlDjCRdj3d
RRRRHIs05CRpRRRRRRRR>R=R
p,RRRRRRRRReRRq pzRRRRRR=>0FF_#H0sM5oRezqp 
2,RRRRRRRRRKRRzQ1aw7Q RR=>Kaz1Q wQ7R,
RRRRRRRRRQRw Rp7RRRR=w>RQ7 p2R;
R8CMRFbsOkC8sFCRI0sHC
;
R-R-R0hFCER0NV0RFmsROD0NR8NMRG]CRNsC8$,RFOkRNMMRF#0R00NsR0IHERRN",3"
-RR-ER0CCRsNH8R#FRVskRMlsLC#FRVs0lN0RC8"Aq3BR"3RCaE#sCRFHk0MRC#o0FRFR
R-0-REMCRCCNs#L0RF8kM##,RFwR"3R "IDHDR0VHR0HMFMRNRH#VGRC858.RF0IMFdR-2R3
RFbsOkC8sBCRE.NsaAsHHR0#5RBRRRRRRRRRRR:RRBRR]qq)B)a ;R
RRRRRRRRRRRRRRRRRRRRRRRRR)z 1pRaRRRRR:kRF0aR17p_zmBtQ_Be a5m).FR8IFM0R;j2
RRRRRRRRRRRRRRRRRRRRRRRRtRRmRm7RRRRR:RRR0FkRmAmph q;R
RRRRRRRRRRRRRRRRRRRRRRRRRQz11 )_ )Rm):MRHRmRAmqp hH2R#R
RLHCoMR
RRNRO#OCRR
H#RRRRRERIC'MRj='R>CRs#0kDRR:=F""j;FRoF:8R=sR0k
C;RRRRRERIC'MR4='R>CRs#0kDRR:=F""4;FRoF:8R=sR0k
C;RRRRRERIC'MR.='R>CRs#0kDRR:=F"".;FRoF:8R=sR0k
C;RRRRRERIC'MRd='R>CRs#0kDRR:=F""d;FRoF:8R=sR0k
C;RRRRRERIC'MRc='R>CRs#0kDRR:=F""c;FRoF:8R=sR0k
C;RRRRRERIC'MR6='R>CRs#0kDRR:=F""6;FRoF:8R=sR0k
C;RRRRRERIC'MRn='R>CRs#0kDRR:=F""n;FRoF:8R=sR0k
C;RRRRRERIC'MR(='R>CRs#0kDRR:=F""(;FRoF:8R=sR0k
C;RRRRRERIC'MRZ='R>CRs#0kDRR:="ZZZ"o;RFRF8:0=Rs;kC
RRRRIRRERCM'RX'=s>RCD#k0=R:RX"XXR";o8FFRR:=0Csk;R
RRRRRIMECREF0CRs#=R>
RRRRRNRR#s#C0FRM01RQ1_z  m)))R
RRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRR"&Rmq) 7sR s:FsRN)C8RRN'&"RR&OR
RRRRRRRR"RR'C,RGObC0RC8NmMROD0NRNOEs0NOC5sRj2-(3R"
RRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRR#sCkRD0:"=Rz"zz;R
RRRRRRFRoFR8RRR:=V#NDCR;
RCRRMO8RN;#C
CRRMb8RsCFO8CksRNBEss.aH0AH#
;
R-R-RsbkbCF#:FR)kM0HCO#RFFllMFR0RC0ER m)qs7RFHk0M
C#RsRbF8OCkRsCmq) 7F_OlMlFRR5
RpRRRRRRRRRRRRRRRRRR:MRHFRk0p Qh;R
RRDR#PRRRRRRRRRRRR:RRR0FkR1RRaz7_pQmtB _eB)am;R
RRoRHFRF8RRRRRRRRR:RRR0FkRARRm mpq
h;RRRRHG8CRRRRRRRRRRRRRF:RkQ0Rhta  
);RRRRO#FM00NMRFLbHRM0:MRHRaQh )t ;RRRRRRR-L-RHsMN$FRbH
M0RRRRO#FM00NMR#lC#CNoRH:RMRRRRmAmph q;R
RRFROMN#0M#0RlEN0R:RRRRHMRARRm mpqRh2H
#
RRRR-b-RkFsb#RC:CFsssCRl#o#NCFRskM0HCR
RRsRbF8OCkRsCClssC5#R
RRRRORRF0M#NRM0l#C#RH:RMaR1)tQh2#RHRRRRRR--CFsssCRl#o#NCR
RRCRLo
HMRRRRRVRHR#lC#CNoRC0EMR
RRRRRRVRHRN#l00ERE
CMRRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRRRRRR"&Rmq) 7V5#H8GC2
R"RRRRRRRRRRRR&CRl#R#
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRCRRD
#CRRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRRRRRR"&Rmq) 7V5kH8GC2
R"RRRRRRRRRRRR&CRl#R#
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRCRRMH8RVR;
RRRRR8CMR;HV
RRRR8CMRFbsOkC8sCCRsCsl#R;
RPRRNNsHLRDCGFoF8RR:Apmm ;qh
RRRRsPNHDNLC$RMLCLDR1:Raz7_pQmtB _eB)amRR5.8MFI0jFR2R;RRRRRR-R-RLdRH
0#RRRRPHNsNCLDR:ORRqB])aqB 
);RRRRPHNsNCLDR:HRRaQh )t ;R
RRNRPsLHNDDCRNk#0RRR:Apmm Rqh:V=RNCD#;RRRRRRR-D-RNR#0OsENNCO0sNRI#MRNR""_
RRRRsPNHDNLCFRVk8M8F:0RRmAmph qRR:=V#NDCR;R-V-RF8kMR8NRF
03RCRLo
HMRRRR1b	H_HIE0bC#NROC5;p2
RRRRRHV#'DPDoCM0>ERR0jRE
CMRRRRRRRH:#=RDEP'H;oE
RRRRsRRCRN85RD,OG,Ro8FF2R;
RRRRRHIEDHCRRj>RRFDFbR
RRRRRRVRHRFGoF=8RRDVN#0CRE
CMRRRRRRRRRsRCs#lCR 5"sssF:MRC8VRFRs#0HRMoCFMOkCM0s"C82R;
RRRRRRRRRHCG0R;
RRRRRCRRDV#HR=ORR''_RC0EMR
RRRRRRRRRHHVRR#=RDDP'C0MoEER0CRM
RRRRRRRRRCRRsCsl#"R5 Fsss1:R0MsHoCRLo#HMR0IHEMRNR_"""2"";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RHVD0N#kER0CRM
RRRRRRRRRCRRsCsl#"R5 Fsssa:RIkFRMs8C#sOFC8#RCO0C0RC8HHMRM0bkRs#0HRMo"_"_"2"";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RC
RRRRRRRRRDRRNk#0RR:=0Csk;R
RRRRRRRRRCRM8H
V;RRRRRRRRCHD#VOR5R'=R3R'20MEC
RRRRRRRRHRRVHR5R4+RRR/=LHbFMR020MEC
RRRRRRRRRRRRsCslRC#5M"COMFk0CCs8"R"3R""NI0RsoFMR8HMC2G";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RHVHRR=#'DPDoCM00ERE
CMRRRRRRRRRRRRClssC5#R"OCMF0kMCN8RR3"""N"R0ER0CCRLoMHMHRMoF0VREDCRH"MC2R;
RRRRRRRRRGRRo8FFRR:=V#NDCR;
RRRRRRRRRCRRG;H0
RRRRRRRRCRRDV#HRkVFMF880ER0CRM
RRRRRRRRRCRRsCsl#"R5aRIF"""3"MRCOMFk0RC8HHMRM0bkRs#0H"Mo2R;
RRRRRRRRRGRRo8FFRR:=V#NDCR;
RRRRRRRRRCRRG;H0
RRRRRRRRCRRMH8RVR;
RRRRRRRRRkVFMF880=R:Rk0sCR;
RRRRRRRRR#DN0:kR=NRVD;#C
RRRRRRRR#CDCR
RRRRRRRRRBsEN.H0sA#H05RO,ML$LDRC,GFoF8l,RCN##o;C2
RRRRRRRRHRRVFRM0oRGFRF80MEC
RRRRRRRRRRRRHCG0R;
RRRRRRRRR8CMR;HV
RRRRRRRR#RRD5PRHFR8IFM0R.H-2=R:RLM$L;DC
RRRRRRRRHRRRR:=HRR-dR;
RRRRRRRRR#DN0:kR=NRVD;#C
RRRRRRRR8CMR;HVRRRRRR
RRRRRRVRHR>HRR0jRE
CMRRRRRRRRRCRsN58RpO,R,oRGF2F8;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRHG8CRR:=HR;
RRRRRFHoF:8R=oRGF;F8
RRRR#CDCR
RRRRRHFoF8=R:Rk0sCR;RRRRRRRRRRRRRRRRR-s-RCRN8HFM0RMNRkRDDNNss$R
RRRRRHG8CRR:=-
4;RRRRCRM8H
V;RMRC8sRbF8OCkRsCmq) 7F_OlMlF;R

RR--hCF0RN0E0FRVsORm0RNDNRM8]RCGs8CN,FR$kNROMFRM00R#NRs0IEH0R"NR3
",R-R-RC0ERNsC8#RHRsVFRlMkL#CsRsVFl0N0C"8RqB3A"R3Ra#ECCFRskM0HCo#RFFR0
-RR-ER0CCRMN#sC0FRLk#M8,FR#R3"w I"RHRDDVRH0HFM0RRNM#GVHC58R.FR8IFM0R2-d3R
RbOsFCs8kC)Rm Rq75RpRR:RRRFHMkp0RQ;h 
RRRRRRRRRRRRRRRRRRRezqp RR:FRk0RhRz)m 1p7e _HkVG2C8R
H#RRRRO#FM00NMRPELRRRR:hRQa  t)=R:R555lHNGl5kld5,Rezqp H'Eo4E+2.2+22/d*-d24R;
RORRF0M#NRM0DRLPR:RRRaQh )t RR:=5H5lMjC5,qRep'z D2FI-/.2dd2*;R
RRNRPsLHND#CRDRPRRRR:1_a7ztpmQeB_ mBa)ER5LDP-L8PRF0IMF2Rj;-RR-HREoLERH
0#RRRRPHNsNCLDRDPNkRCG:hRz)m 1p7e _HkVGRC85PELRI8FMR0FD2LP;R
RRNRPsLHNDHCRo8FFRRR:Apmm ;qh
RRRRsPNHDNLCRRHRRRRRQ:Rhta  
);RCRLo
HMRRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;
RmRR)7 q_lOFlRFM5RRp=p>R,R
RRRRRRRRRRRRRRRRRRP#DRR=>#,DP
RRRRRRRRRRRRRRRRRRRHFoF8>R=RFHoF
8,RRRRRRRRRRRRRRRRRHRR8RCG=H>R,R
RRRRRRRRRRRRRRRRRRFLbHRM0=->RD,LP
RRRRRRRRRRRRRRRRRRRl#C#NRoC=0>Rs,kC
RRRRRRRRRRRRRRRRRRR#0lNE>R=RDVN#;C2
RRRRRHVHFoF8ER0CRMRRRRRRRRRRRRRRRRRRRRRRR--W8CRHM8RFo0RCN0RMEF0CCsRsssF
RRRRHRRVFRM05R5HRR=-R42NRM8RRRRRRRRRRRRR-R-RRWCs8CNRCCPsE$0H,MoR8NMRoEHEHRL0j#R
RRRRRRRRRRRR5RRF5sR#5DPE-LPDRLP8MFI0eFRq pz'oEHE-+4D2LP2RR='2j'2ER0CRM
RRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRRR&mR")7 q5HkVG2C8:CReOs0FRk0sM0ONC"83
RRRRRRRR#RRCsPCHR0$CFsssR;
RRRRR#CDCR
RRRRRRVRHRs5FRD5#Pq5ep'z D-FID-LP4FR8IFM0R2j2R'=R4R'20MEC
RRRRRRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRRRRRR&mR")7 q5HkVG2C8:CReOs0FRk0sM0ONC
8"RRRRRRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRRMRC8VRH;R
RRRRRRNRPDGkCRR:=0kF_VCHG8#R5DRP,E,LPRPDL2R;
RRRRReRRq pzR=R:RDPNkRCG5peqzs 'NCMo2R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMb8RsCFO8CksR m)q
7;
bRRsCFO8CksR m)qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_kH8GC;R
RRRRRRRRRRRRRRRRRt7mmRRR:FRk0RmRAmqp hH2R#R
RRFROMN#0ME0RLRPRRRR:Q hatR ):5=R5N5lGkHll,5dRq5ep'z EEHo+242+/.2dd2*2;-4
RRRRMOF#M0N0LRDPRRRRQ:Rhta  :)R=5R5lCHM5Rj,ezqp F'DI.2-22/d*
d;RRRRPHNsNCLDRP#DRRRR:aR17p_zmBtQ_Be aRm)5PEL-PDLRI8FMR0FjR2;RR--EEHoR0LH#R
RRNRPsLHNDPCRNCDkGRR:z h)1emp k7_VCHG8ER5L8PRF0IMFLRDP
2;RRRRPHNsNCLDRFHoFR8R:mRAmqp hR;
RPRRNNsHLRDCHRRRR:RRRaQh )t ;R
RLHCoMR
RRqRepRz :5=Rezqp N'sMRoC='>Rz;'2
RRRR m)qO7_FFllMRR5p>R=R
p,RRRRRRRRRRRRRRRRR#RRD=PR>DR#PR,
RRRRRRRRRRRRRRRRRoRHFRF8=H>Ro8FF,R
RRRRRRRRRRRRRRRRRRCH8G>R=R
H,RRRRRRRRRRRRRRRRRLRRbMFH0>R=RL-DPR,
RRRRRRRRRRRRRRRRRCRl#o#NC>R=RDVN#
C,RRRRRRRRRRRRRRRRR#RRlEN0RR=>V#NDC
2;RRRRH5VRHFoF8MRN8RRRRRRRRRRRRRRRRRRR-W-RCHR88FRM0CRo0MRNFC0EssRCs
FsRRRRRRRR5=HRR2-4R8NMRRRRRRRRRRRRRRRR-W-RCCRsNC8RP$Cs0MEHoN,RME8RHRoEL#H0RRj
RRRRR5RRF5sR#5DPE-LPDRLP8MFI0eFRq pz'oEHE-+4D2LP2RR='2j'2ER0CRM
RRRRRDPNkRCG:0=RFV_kH8GCRD5#PE,RLRP,D2LP;R
RRRRRezqp :RR=NRPDGkCRq5ep'z soNMC
2;RRRRRFRoF:8R=sR0k
C;RRRRCCD#
RRRRoRRFRF8:V=RNCD#;R
RRMRC8VRH;R
RCRM8bOsFCs8kC)Rm ;q7
R
RbOsFCs8kC)Rm 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp #7_VCHG8H2R#R
RRFROMN#0ME0RLRPRRRR:Q hatR ):5=R5N5lGkHll,5dRq5ep'z EEHo+242+/.2dd2*2;-4
RRRRMOF#M0N0LRDPRRRRQ:Rhta  :)R=5R5lCHM5Rj,ezqp F'DI.2-22/d*
d;RRRRPHNsNCLDRP#DRRRR:aR17p_zmBtQ_Be aRm)5PEL-PDLRI8FMR0FjR2;RR--EEHoR0LH#R
RRNRPsLHNDPCRNCDkGRR:z h)1emp #7_VCHG8ER5L8PRF0IMFLRDP
2;RRRRPHNsNCLDRFHoFR8R:mRAmqp hR;
RPRRNNsHLRDCHRRRR:RRRaQh )t ;R
RLHCoMR
RRqRepRz :5=Rezqp N'sMRoC='>Rz;'2
RRRR m)qO7_FFllMRR5p>R=R
p,RRRRRRRRRRRRRRRRR#RRD=PR>DR#PR,
RRRRRRRRRRRRRRRRRoRHFRF8=H>Ro8FF,R
RRRRRRRRRRRRRRRRRRCH8G>R=R
H,RRRRRRRRRRRRRRRRRLRRbMFH0>R=RL-DPR,
RRRRRRRRRRRRRRRRRCRl#o#NC>R=Rk0sCR,
RRRRRRRRRRRRRRRRRlR#NR0E=0>Rs2kC;R
RRVRHRFHoF08RERCMRRRRRRRRRRRRRRRRRRRRR-R-RRWC8RH8MRF0oRC0N0MFERCsCFsssR
RRRRRHMVRF50R5=HRR2-4R8NMRRRRRRRRRRRRR-RR-CRWRNsC8PRCC0s$EoHM
RRRRRRRRRRRR5RR5P#D5peqzE 'H-oED2LPR'=RjN'RMR8RRRRR-#-RHRoML#H0RC=RGN0sR0LH#R
RRRRRRRRRRRRRRsRFRD5#PL5EPL-DPFR8IFM0RpeqzE 'H+oE4L-DPR22=jR''F2RsR
RRRRRRRRRRRRRRD5#Pq5ep'z EEHo-PDL2RR='R4'N
M8RRRRRRRRRRRRRRRRNRM85P#D5PEL-PDLRI8FMR0Fezqp H'Eo4E+-PDL2=2RR''42R220MEC
RRRRRRRRbsCFRs0VCHG8	_boM'H#M0NOMC_N
lCRRRRRRRRRRR&" m)q#75VCHG8R2:e0COF0sRsOkMN80C3R"
RRRRRRRRRP#CC0sH$sRCs;Fs
RRRRCRRD
#CRRRRRRRRH5VRF5sR#5DPezqp F'DIL-DPR-48MFI0jFR2=2RR''42ER0CRM
RRRRRRRRR#N#CRs0hWm_qQ)hhRt
RRRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRRRRRR&" m)q#75VCHG8R2:e0COF0sRsOkMN80C"R
RRRRRRRRRRCR#PHCs0I$RNHsMM
o;RRRRRRRRCRM8H
V;RRRRRRRRPkNDC:GR=FR0_H#VGRC85P#D,LREPD,RL;P2
RRRRRRRRpeqzR R:P=RNCDkGeR5q pz'MsNo;C2
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRFbsOkC8smCR)7 q;R

RFbsOkC8smCR)7 q5RpRR:RRRFHMkp0RQ;h 
RRRRRRRRRRRRRRRReRRq pzRF:RkR0RR)zh p1me_ 7#GVHC
8;RRRRRRRRRRRRRRRRRmRtmR7R:kRF0RRRApmm 2qhR
H#RRRRO#FM00NMRPELRRRR:hRQa  t)=R:R555lHNGl5kld5,Rezqp H'Eo4E+2.2+22/d*-d24R;
RORRF0M#NRM0DRLPR:RRRaQh )t RR:=5H5lMjC5,qRep'z D2FI-/.2dd2*;R
RRNRPsLHND#CRDRPRRRR:1_a7ztpmQeB_ mBa)ER5LDP-L8PRF0IMF2Rj;-RR-HREoLERH
0#RRRRPHNsNCLDRDPNkRCG:hRz)m 1p7e _H#VGRC85PELRI8FMR0FD2LP;R
RRNRPsLHNDHCRo8FFRRR:Apmm ;qh
RRRRsPNHDNLCRRHRRRRRQ:Rhta  
);RCRLo
HMRRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;
RmRR)7 q_lOFlRFM5RRp=p>R,R
RRRRRRRRRRRRRRRRRRP#DRR=>#,DP
RRRRRRRRRRRRRRRRRRRHFoF8>R=RFHoF
8,RRRRRRRRRRRRRRRRRHRR8RCG=H>R,R
RRRRRRRRRRRRRRRRRRFLbHRM0=->RD,LP
RRRRRRRRRRRRRRRRRRRl#C#NRoC=V>RNCD#,R
RRRRRRRRRRRRRRRRRRN#l0=ER>sR0k;C2
RRRRRHV5FHoFR8RRRRRRRRRRRRRRRRRRRRRRR--W8CRHM8RFo0RCN0RMEF0CCsRsssF
RRRRRRRR8NMRR5H=4R-2RRRRRRRRRRRRRRRRR--WsCRCRN8CsPC$H0EMRo
RRRRRNRRM58R5P#D5peqzE 'H-oED2LPR'=RjN'RMR8R-#-RHRoML#H0RC=RGN0sR0LH#R
RRRRRRRRRRRRRF5sR#5DPE-LPDRLP8MFI0eFRq pz'oEHE-+4D2LP2RR='2j'R
FsRRRRRRRRRRRRRD5#Pq5ep'z EEHo-PDL2RR='R4'N
M8RRRRRRRRRRRRRMRN8#R5DEP5LDP-L8PRF0IMFqRep'z EEHo+D4-L2P2R'=R42'22ER0CRM
RRRRRDPNkRCG:0=RFV_#H8GCRD5#PE,RLRP,D2LP;R
RRRRRezqp :RR=NRPDGkCRq5ep'z soNMC
2;RRRRRFRoF:8R=sR0k
C;RRRRCCD#
RRRRoRRFRF8:V=RNCD#;R
RRMRC8VRH;R
RCRM8bOsFCs8kC)Rm ;q7
R
R-E-RCsGRCRN8NRM8I0sHCR
RbOsFCs8kCIREsCH0RR5
RpRRRRRRRRRRRH:RM0FkRhpQ R;RRRRRRRRRRRRRRR--HkMb0HRDMRC
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7kGVHCR8;RR--VCHG8FRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RH
LRRCMoHR-R-RN GlCbDR3jddRj
RIRRsCH0RR5pRRRRRRRR=p>R,R
RRRRRRRRRRpeqzR RR=RR>FR0_0E#soHMRq5ep2z ,R
RRRRRRRRRR1KzaQQw =7R>zRK1waQQ, 7
RRRRRRRRRRRwpQ 7RRRR>R=R wQp;72
CRRMb8RsCFO8CksRsEIH;0C
R
R-b-RkFsb#RC:I0sHCV#RH8GCRHbFMH0RMR0FNHRDMRC
RFbsOkC8sECRI0sHC
R5RRRRpRRRRRRRRRR:HkMF0QRphR ;RRRRRRRRRRRRR-R-RbHMkD0RH
MCRRRRezqp RRRRRR:HRMRRhRz)m 1p7e _H#VG;C8R-R-RGVHCb8RF0HMRbHMkR0
RKRRzQ1aw7Q RH:RMRRRR71Q :RR=HRso;E0
RRRR wQpR7RR:RRRRHMRWRRQ]7aRR:=jH2R#R
RLHCoM-RR-GR NDlbCdRj3
djRRRRI0sHCpR5RRRRRRRRRR=>pR,
RRRRRRRRRqRepRz RRRR=0>RF#_E0MsHoeR5q pz2R,
RRRRRRRRRzRK1waQQR 7=K>RzQ1aw7Q ,R
RRRRRRRRRR wQpR7RR=RR>QRw 2p7;R
RCRM8bOsFCs8kCIREsCH0;R

RR--]RCG)8CNR8NMRHWs0bCRsCFO8Cks#FRVsaR17p_zmBtQ_Be a3m)
-RR-FRv8HHVCV8RsRFl0RECFosHHDMNRR0FLlCRFRsCVoFsHMPHo
3
RsRbF8OCkRsCBsEN.NTk80AH#BR5RRRRRRRRR:RRRRRRRqB])aqB 
);RRRRRRRRRRRRRRRRRRRRRRRRR)RR p1zaRRRR:RRR0FkR71a_mzpt_QBea Bmd)5RI8FMR0Fj
2;RRRRRRRRRRRRRRRRRRRRRRRRRtRRmRm7RRRRR:RRR0FkRmAmph q;R
RRRRRRRRRRRRRRRRRRRRRRRRRR1Q1z  _)))mRH:RMARRm mpqRh2HR#
RoLCHRM
RORRNR#CO#RH
RRRRIRRERCM'Rj'RRRRR>R=R#sCkRD0:G=R";j"RFoF8=R:Rk0sCR;
RRRRRCIEM4R''RRRRRRR=s>RCD#k0=R:R4G""o;RFRF8:0=Rs;kC
RRRRIRRERCM'R.'RRRRR>R=R#sCkRD0:G=R";."RFoF8=R:Rk0sCR;
RRRRRCIEMdR''RRRRRRR=s>RCD#k0=R:RdG""o;RFRF8:0=Rs;kC
RRRRIRRERCM'Rc'RRRRR>R=R#sCkRD0:G=R";c"RFoF8=R:Rk0sCR;
RRRRRCIEM6R''RRRRRRR=s>RCD#k0=R:R6G""o;RFRF8:0=Rs;kC
RRRRIRRERCM'Rn'RRRRR>R=R#sCkRD0:G=R";n"RFoF8=R:Rk0sCR;
RRRRRCIEM(R''RRRRRRR=s>RCD#k0=R:R(G""o;RFRF8:0=Rs;kC
RRRRIRRERCM'RU'RRRRR>R=R#sCkRD0:G=R";U"RFoF8=R:Rk0sCR;
RRRRRCIEMgR''RRRRRRR=s>RCD#k0=R:RgG""o;RFRF8:0=Rs;kC
RRRRIRRERCM'Rq'|NR''>R=R#sCkRD0:G=R";q"RFoF8=R:Rk0sCR;
RRRRRCIEMAR''RR|'RL'=s>RCD#k0=R:RAG""o;RFRF8:0=Rs;kC
RRRRIRRERCM'RB'|OR''>R=R#sCkRD0:G=R";B"RFoF8=R:Rk0sCR;
RRRRRCIEM7R''RR|'R8'=s>RCD#k0=R:R7G""o;RFRF8:0=Rs;kC
RRRRIRRERCM'R '|CR''>R=R#sCkRD0:G=R"; "RFoF8=R:Rk0sCR;
RRRRRCIEMwR''RR|'RV'=s>RCD#k0=R:RwG""o;RFRF8:0=Rs;kC
RRRRIRRERCM'RZ'RRRRR>R=R#sCkRD0:"=RZZZZ"o;RFRF8:0=Rs;kC
RRRRIRRERCM'RX'RRRRR>R=R#sCkRD0:"=RXXXX"o;RFRF8:0=Rs;kC
RRRRIRRERCMFC0Es=#R>R
RRRRRR#RN#0CsR0MFR1Q1z  _)))m
RRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRRR&]R")7 qRs sFRs:)8CNR'NR"RR&O
R&RRRRRRRRR'R",GRCb0COCN8RRG]CRNOEs0NOC5sRj2-w3R"
RRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRR#sCkRD0:"=Rzzzz"R;
RRRRRoRRFRF8R=R:RDVN#
C;RRRRCRM8OCN#;R
RCRM8bOsFCs8kCERBNTs.kAN8H;0#
R
R-b-RkFsb#RC:)0FkH#MCRlOFlRFM00FRE]CR)7 qRksF0CHM#R
RbOsFCs8kC)R] _q7OlFlF5MR
RRRRRpRRRRRRRRRRRRRRRR:HkMF0QRph
 ;RRRR#RDPRRRRRRRRRRRRRF:RkR0RR71a_mzpt_QBea Bm
);RRRRHFoF8RRRRRRRRRRRRF:RkR0RRmAmph q;R
RR8RHCRGRRRRRRRRRR:RRR0FkRaQh )t ;R
RRFROMN#0ML0RbMFH0RR:HQMRhta  R);RRRRR-R-RMLHNRs$bMFH0R
RRFROMN#0Ml0RCN##o:CRRRHMRARRm mpq
h;RRRRO#FM00NMRN#l0RERRH:RMRRRRmAmph q2#RH
R
RR-R-RsbkbCF#:sRCsRFsl#C#NRoCs0FkH
MCRRRRbOsFCs8kCsRCs#lCRR5
RRRRRMOF#M0N0CRl#:#RRRHM1Qa)hRt2HR#RR-RR-sRCsRFsl#C#N
oCRRRRLHCoMR
RRRRRHlVRCN##o0CRE
CMRRRRRRRRH#VRlEN0RC0EMR
RRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRR&RRR)"] 5q7#GVHCR82"R
RRRRRRRRRRRR&l#C#
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRR#CDCR
RRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRR&RRR)"] 5q7kGVHCR82"R
RRRRRRRRRRRR&l#C#
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RCRRMb8RsCFO8CksRsCsl;C#
RRRRsPNHDNLCoRGFRF8RA:Rm mpq
h;RRRRPHNsNCLDRLM$LRDC:aR17p_zmBtQ_Be aRm)58dRF0IMF2Rj;RRRRRRRRR--cHRL0R#
RPRRNNsHLRDCORRRR:RRRqB])aqB 
);RRRRPHNsNCLDRRHRRRRR:hRQa  t)R;
RPRRNNsHLRDCD0N#k:RRRmAmph qRR:=V#NDCR;RRRRRRR--D0N#RNOEs0NOCIsRNN#RM_R""R
RRNRPsLHNDVCRF8kM8RF0:mRAmqp h=R:RDVN#RC;RR--VMFk8RRN83F0
LRRCMoH
RRRRH1	bE_IH#0CbCNOR25p;RRR
RRRRRHV#'DPDoCM0>ERR0jRE
CMRRRRRRRH:#=RDEP'H;oE
RRRRsRRCRN85RD,OG,Ro8FF2R;
RRRRRHIEDHCRRj>RRFDFbR
RRRRRRVRHRFGoF=8RRDVN#0CRE
CMRRRRRRRRRsRCs#lCR 5"sssF:MRC8VRFRs#0HRMoCFMOkCM0s"C82R;
RRRRRRRRRHCG0R;
RRRRRCRRDV#HR=ORR''_RC0EMR
RRRRRRRRRHHVRR#=RDDP'C0MoEER0CRM
RRRRRRRRRCRRsCsl#"R5 Fsss1:R0MsHoCRLo#HMR0IHEMRNR_"""2"";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RHVD0N#kER0CRM
RRRRRRRRRCRRsCsl#"R5 Fsssa:RIkFRMs8C#sOFC8#RCO0C0RC8HHMRM0bkRs#0HRMo"_"_"2"";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RC
RRRRRRRRRDRRNk#0RR:=0Csk;R
RRRRRRRRRCRM8H
V;RRRRRRRRCHD#VOR5R'=R3R'20MEC
RRRRRRRRHRRVHR5R4+RRR/=LHbFMR020MEC
RRRRRRRRRRRRsCslRC#5M"COMFk0CCs8"R"3R""NI0RsoFMR8HMC2G";R
RRRRRRRRRRoRGFRF8:V=RNCD#;R
RRRRRRRRRRGRCH
0;RRRRRRRRRDRC#RHVHRR=#'DPDoCM00ERE
CMRRRRRRRRRRRRClssC5#R"OCMF0kMCN8RR3"""N"R0ER0CCRLoMHMHRMoF0VREDCRH"MC2R;
RRRRRRRRRGRRo8FFRR:=V#NDCR;
RRRRRRRRRCRRG;H0
RRRRRRRRCRRDV#HRkVFMF880ER0CRM
RRRRRRRRRCRRsCsl#"R5aRIF"""3"MRCOMFk0RC8HHMRM0bkRs#0H"Mo2R;
RRRRRRRRRGRRo8FFRR:=V#NDCR;
RRRRRRRRRCRRG;H0
RRRRRRRRCRRMH8RVR;
RRRRRRRRRkVFMF880=R:Rk0sCR;
RRRRRRRRR#DN0:kR=NRVD;#C
RRRRRRRR#CDCR
RRRRRRRRRBsEN.NTk80AH#,5ORLM$L,DCRFGoFR8,l#C#N2oC;R
RRRRRRRRRHMVRFG0Ro8FFRC0EMR
RRRRRRRRRRGRCH
0;RRRRRRRRRMRC8VRH;R
RRRRRRRRR#RDP58HRF0IMF-RHd:2R=$RMLCLD;R
RRRRRRRRRH=R:R-HRR
c;RRRRRRRRRNRD#R0k:V=RNCD#;R
RRRRRRMRC8VRH;RRRRRR
RRRRRHRRVRRH>RRj0MEC
RRRRRRRRsRRCRN85Rp,OG,Ro8FF2R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRCH8G=R:R
H;RRRRRoRHFRF8:G=Ro8FF;R
RRDRC#RC
RRRRRCH8G=R:R;-4
RRRRHRRo8FFRR:=0Csk;RRRRRRRRRRRRRRRRRRRRR--s8CNRDMkD0R#soHM
RRRR8CMR;HV
CRRMb8RsCFO8CksR ])qO7_FFllM
;
RsRbF8OCkRsC]q) 7R5pRRRR:MRHFRk0p Qh;R
RRRRRRRRRRRRRRRRRezqp RR:FRk0RhRz)m 1p7e _HkVG2C8R
H#RRRRO#FM00NMRPELRRRR:hRQa  t)=R:R555lHNGl5klc5,Rezqp H'Eo4E+2d2+22/c*-c24R;
RORRF0M#NRM0DRLPR:RRRaQh )t RR:=5H5lMjC5,qRep'z D2FI-/d2cc2*;R
RRNRPsLHND#CRDRPRRRR:1_a7ztpmQeB_ mBa)ER5LDP-L8PRF0IMF2Rj;-RR-HREoLERH
0#RRRRPHNsNCLDRDPNkRCG:hRz)m 1p7e _HkVGRC85PELRI8FMR0FD2LP;R
RRNRPsLHNDHCRo8FFRRR:Apmm ;qh
RRRRsPNHDNLCRRHRRRRRQ:Rhta  
);RCRLo
HMRRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;
R]RR)7 q_lOFlRFM5RRp=p>R,R
RRRRRRRRRRRRRRRRRRP#DRR=>#,DP
RRRRRRRRRRRRRRRRRRRHFoF8>R=RFHoF
8,RRRRRRRRRRRRRRRRRHRR8RCG=H>R,R
RRRRRRRRRRRRRRRRRRFLbHRM0=->RD,LP
RRRRRRRRRRRRRRRRRRRl#C#NRoC=V>RNCD#,R
RRRRRRRRRRRRRRRRRRN#l0=ER>NRVD2#C;R
RRVRHRFHoF08RE
CMRRRRRVRHR0MFRH55R-=R4N2RMR8RRRRRRRRRRRRRRR--WsCRCRN8CsPC$H0EMRo,NRM8EEHoR0LH#
RjRRRRRRRRRRRRRFR5s#R5DEP5LDP-L8PRF0IMFqRep'z EEHo+D4-L2P2R'=Rj2'2RC0EMR
RRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRR&RRR)"] 5q7kGVHC:82ROeC0RFs0MskOCN08
3"RRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRCCD#
RRRRRRRRRHV5RFs5P#D5peqzD 'FDI-L4P-RI8FMR0FjR22=4R''02RE
CMRRRRRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRR&RRR)"] 5q7kGVHC:82ROeC0RFs0MskOCN08R"
RRRRRRRRR#RRCsPCHR0$IMNsH;Mo
RRRRRRRR8CMR;HV
RRRRRRRRDPNkRCG:0=RFV_kH8GCRD5#PE,RLRP,D2LP;R
RRRRRRqRepRz RR:=PkNDC5GRezqp N'sM2oC;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8sRbF8OCkRsC]q) 7
;
RsRbF8OCkRsC]q) 7R5pRRRR:MRHFRk0p Qh;R
RRRRRRRRRRRRRRRRRezqp RR:FRk0RhRz)m 1p7e _HkVG;C8
RRRRRRRRRRRRRRRRtRRmRm7RF:RkR0RRmAmph q2#RH
RRRRMOF#M0N0LREPRRRRQ:Rhta  :)R=5R55GlNHllk5Rc,5peqzE 'H+oE4+22dc2/22*c-
4;RRRRO#FM00NMRPDLRRRR:hRQa  t)=R:Rl55H5MCje,Rq pz'IDF22-d/*c2cR;
RPRRNNsHLRDC#RDPR:RRR71a_mzpt_QBea Bm5)RE-LPDRLP8MFI0jFR2R;R-E-RHRoEL#H0
RRRRsPNHDNLCNRPDGkCRz:Rh1) m pe7V_kH8GCRL5EPFR8IFM0RPDL2R;
RPRRNNsHLRDCHFoF8:RRRmAmph q;R
RRNRPsLHNDHCRRRRRRRR:Q hat; )
LRRCMoH
RRRRpeqz: R=eR5q pz'MsNo=CR>zR''
2;RRRR]q) 7F_OlMlFRp5RRR=>pR,
RRRRRRRRRRRRRRRRRDR#P>R=RP#D,R
RRRRRRRRRRRRRRRRRRFHoF=8R>oRHF,F8
RRRRRRRRRRRRRRRRRRRHG8CRR=>HR,
RRRRRRRRRRRRRRRRRbRLF0HMRR=>-PDL,R
RRRRRRRRRRRRRRRRRR#lC#CNoRR=>V#NDCR,
RRRRRRRRRRRRRRRRRlR#NR0E=V>RNCD#2R;
RHRRVHR5o8FFR8NMRRRRRRRRRRRRRRRRR-RR-CRWR88HR0MFR0oCRFNM0sECRsCsFRs
RRRRR5RRHRR=-R42NRM8RRRRRRRRRRRRR-RR-CRWRNsC8PRCC0s$EoHM,MRN8HREoLERHR0#jR
RRRRRRFR5s#R5DEP5LDP-L8PRF0IMFqRep'z EEHo+D4-L2P2R'=Rj2'2RC0EMR
RRRRRPkNDC:GR=FR0_HkVGRC85P#D,LREPD,RL;P2
RRRReRRq pzR=R:RDPNkRCG5peqzs 'NCMo2R;
RRRRRFoF8=R:Rk0sCR;
RCRRD
#CRRRRRFRoF:8R=NRVD;#C
RRRR8CMR;HV
CRRMb8RsCFO8CksR ])q
7;
bRRsCFO8CksR ])qp75RRRRRH:RM0FkRhpQ R;
RRRRRRRRRRRRRRRRRpeqz: RR0FkRzRRh1) m pe7V_#H8GC2#RH
RRRRMOF#M0N0LREPRRRRQ:Rhta  :)R=5R55GlNHllk5Rc,5peqzE 'H+oE4+22dc2/22*c-
4;RRRRO#FM00NMRPDLRRRR:hRQa  t)=R:Rl55H5MCje,Rq pz'IDF22-d/*c2cR;
RPRRNNsHLRDC#RDPR:RRR71a_mzpt_QBea Bm5)RE-LPDRLP8MFI0jFR2R;R-E-RHRoEL#H0
RRRRsPNHDNLCNRPDGkCRz:Rh1) m pe7V_#H8GCRL5EPFR8IFM0RPDL2R;
RPRRNNsHLRDCHFoF8:RRRmAmph q;R
RRNRPsLHNDHCRRRRRRRR:Q hat; )
LRRCMoH
RRRRpeqz: R=eR5q pz'MsNo=CR>zR''
2;RRRR]q) 7F_OlMlFRp5RRR=>pR,
RRRRRRRRRRRRRRRRRDR#P>R=RP#D,R
RRRRRRRRRRRRRRRRRRFHoF=8R>oRHF,F8
RRRRRRRRRRRRRRRRRRRHG8CRR=>HR,
RRRRRRRRRRRRRRRRRbRLF0HMRR=>-PDL,R
RRRRRRRRRRRRRRRRRR#lC#CNoRR=>0Csk,R
RRRRRRRRRRRRRRRRRRN#l0=ER>sR0k;C2
RRRRRHVHFoF8ER0CRMRRRRRRRRRRRRRRRRRRRRRRR--W8CRHM8RFo0RCN0RMEF0CCsRsssF
RRRRHRRVFRM05R5HRR=-R42RRRRRRRRRRRRRRRRR-R-RRWCs8CNRCCPsE$0H
MoRRRRRRRRRRRRRMRN85R5#5DPezqp H'EoDE-LRP2=jR''MRN8-RR-HR#oLMRHR0#=GRC0RsNL#H0
RRRRRRRRRRRRRRRRRRRRRFs5P#D5PEL-PDLRI8FMR0Fezqp H'Eo4E+-PDL2=2RR''j2sRF
RRRRRRRRRRRRRRRRRRR5P#D5peqzE 'H-oED2LPR'=R4N'RMR8
RRRRRRRRRRRRRRRRRNRRM58R#5DPE-LPDRLP8MFI0eFRq pz'oEHE-+4D2LP2RR='24'202RE
CMRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRR"&R]q) 7V5#H8GC2e:RCFO0ssR0kNMO03C8"R
RRRRRRRRR#CCPs$H0RsCsF
s;RRRRRDRC#RC
RRRRRHRRVFR5s#R5DeP5q pz'IDF-PDL-84RF0IMF2Rj2RR='24'RC0EMR
RRRRRRRRRNC##sh0Rmq_W)hhQtR
RRRRRRRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRRRRRRRRRR"&R]q) 7V5#H8GC2e:RCFO0ssR0kNMO0"C8
RRRRRRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRRCRRMH8RVR;
RRRRRPRRNCDkG=R:R_0F#GVHC58R#,DPRPEL,LRDP
2;RRRRRRRRezqp :RR=NRPDGkCRq5ep'z soNMC
2;RRRRRMRC8VRH;R
RRMRC8VRH;R
RCRM8bOsFCs8kC)R] ;q7
R
RbOsFCs8kC)R] 5q7pRRRRRR:HkMF0QRph
 ;RRRRRRRRRRRRRRRRRqRepRz :kRF0RRRz h)1emp #7_VCHG8R;
RRRRRRRRRRRRRRRRRmtm7:RRR0FkRARRm mpqRh2HR#
RORRF0M#NRM0ERLPR:RRRaQh )t RR:=5l55NlGHkcl5,eR5q pz'oEHE2+422+d/*c2c42-;R
RRFROMN#0MD0RLRPRRRR:Q hatR ):5=R5MlHC,5jRpeqzD 'F-I2dc2/2;*c
RRRRsPNHDNLCDR#PRRRR1:Raz7_pQmtB _eB)amRL5EPL-DPFR8IFM0R;j2R-R-RoEHEHRL0R#
RPRRNNsHLRDCPkNDC:GRR)zh p1me_ 7#GVHC58RERLP8MFI0DFRL;P2
RRRRsPNHDNLCoRHFRF8RA:Rm mpq
h;RRRRPHNsNCLDRRHRRRRR:hRQa  t)R;
RoLCHRM
ReRRq pzRR:=5peqzs 'NCMoRR=>'2z';R
RR)R] _q7OlFlF5MRR=pR>,Rp
RRRRRRRRRRRRRRRRRRR#RDP=#>RD
P,RRRRRRRRRRRRRRRRRHRRo8FFRR=>HFoF8R,
RRRRRRRRRRRRRRRRR8RHC=GR>,RH
RRRRRRRRRRRRRRRRRRRLHbFM=0R>DR-L
P,RRRRRRRRRRRRRRRRRlRRCN##o=CR>NRVD,#C
RRRRRRRRRRRRRRRRRRR#0lNE>R=Rk0sC
2;RRRRH5VRHFoF8MRN8RRRRRRRRRRRRRRRRRRR-W-RCHR88FRM0CRo0MRNFC0EssRCs
FsRRRRRRRR5=HRR2-4R8NMRRRRRRRRRRRRRRRR-W-RCCRsNC8RP$Cs0MEHoR
RRRRRR5R5#5DPezqp H'EoDE-LRP2=jR''MRN8-RR-HR#oLMRHR0#=GRC0RsNL#H0
RRRRRRRRFRRs#R5DEP5LDP-L8PRF0IMFqRep'z EEHo+D4-L2P2R'=RjR'2FRs
RRRRRRRR5P#D5peqzE 'H-oED2LPR'=R4N'RMR8
RRRRRRRRR8NMRD5#PL5EPL-DPFR8IFM0RpeqzE 'H+oE4L-DPR22=4R''222RC0EMR
RRRRRPkNDC:GR=FR0_H#VGRC85P#D,LREPD,RL;P2
RRRReRRq pzR=R:RDPNkRCG5peqzs 'NCMo2R;
RRRRRFoF8=R:Rk0sCR;
RCRRD
#CRRRRRFRoF:8R=NRVD;#C
RRRR8CMR;HV
CRRMb8RsCFO8CksR ])q
7;
-RR-FRa_s#0HRMoVOkM0MHF#R3RzV#CkHDRMsR"CsbF0#"R0CN0l0CM#R3
RR-- lGNb:DCRCRsb0FsRC"s#0kDR#INR&"RR_0F#H0sMso5CD#k0
2;RkRVMHO0F0MRF0_#soHMRN5PDRkC:hRz)m 1p7e _HkVG2C8R0sCkRsM1Qa)hHtR#R
RRNRPsLHND#CRRRRRR1:Rah)QtR540PFRNCDk'MDCoR0E+R42:5=RFC0Es=#R>RR''
2;RRRRPHNsNCLDRL#kPRND:hRz)m 1p7e _HkVGRC85DPNkEC'HRoE8MFI0-FR4
2;RRRRPHNsNCLDRM#H8:GRRaQh )t ;R
RLHCoMR
RRVRHRDPNkDC'C0MoERR<4ER0CRM
RRRRR0sCkRsMh;z1
RRRR#CDCR
RRRRRHPVRNCDk'oEHERR<jER0CRM
RRRRRHRRVNRPD5kCPkNDCH'EoRE2=ZR''ER0CRM
RRRRRRRRR0sCkRsM0#F_0MsHosR5Cx#HC#R5VCHG8N5PD2kC,,RjRDPNkDC'F2I2;R
RRRRRRDRC#RC
RRRRRRRRR0sCkRsM0#F_0MsHosR5Cx#HCPR5NCDk,,RjRDPNkDC'F2I2;R
RRRRRRMRC8VRH;R
RRRRRCHD#VNRPD'kCDRFI>j=RRC0EMR
RRRRRRVRHR_Q#XPR5NCDk5DPNkDC'F2I2RC0EMR
RRRRRRRRR#PkLN:DR=FR50sEC#>R=RDPNkPC5NCDk'IDF2
2;RRRRRRRRRkR#LDPNRN5PD'kCsoNMC:2R=NRPD;kC
RRRRRRRRsRRCs0kMFR0_s#0H5Mo#PkLN;D2
RRRRRRRR#CDCR
RRRRRRRRRskC0s0MRF0_#soHMRC5s#CHxRN5PD,kCRDPNkEC'H,oER2-42R;
RRRRRCRRMH8RVR;
RRRRR#CDCR
RRRRRRHR#MR8G:4=R;R
RRRRRRFRVsRRHHPMRNCDk'oEHEFR8IFM0RDPNkDC'FDIRF
FbRRRRRRRRRVRHR=HRRR-40MEC
RRRRRRRRRRRR##5HGM82=R:R''3;R
RRRRRRRRRRHR#MR8GR:RR=HR#MR8G+;R4
RRRRRRRRCRRMH8RVR;
RRRRRRRRR##5HGM82=R:RpvegF_0_NOEsa517p_zmBtQ5DPNkHC52;22
RRRRRRRR#RRHGM8RRRR:#=RHGM8R4+R;R
RRRRRRMRC8FRDF
b;RRRRRRRRskC0s#MR;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F0MRF0_#soHM;R

RMVkOF0HMFR0_s#0HRMo5DPNk:CRR)zh p1me_ 7#GVHCR82skC0s1MRah)Qt#RH
RRRRsPNHDNLCRR#RRRR:aR1)tQh504RFNRPD'kCDoCM0+ERRR42:5=RFC0Es=#R>RR''
2;RRRRPHNsNCLDRL#kPRND:hRz)m 1p7e _H#VGRC85DPNkEC'HRoE8MFI0-FR4
2;RRRRPHNsNCLDRM#H8:GRRaQh )t ;R
RLHCoMR
RRVRHRDPNkDC'C0MoERR<4ER0CRM
RRRRR0sCkRsMh;z1
RRRR#CDCR
RRRRRHPVRNCDk'oEHERR<jER0CRM
RRRRRsRRCs0kMFR0_s#0HRMo5#sCHRxC5DPNkRC,jP,RNCDk'IDF2
2;RRRRRDRC#RHVPkNDCF'DI=R>R0jRE
CMRRRRRRRRHQVR#R_X5DPNkPC5NCDk'IDF202RE
CMRRRRRRRRRkR#LDPNRR:=5EF0CRs#=P>RNCDk5DPNkDC'F2I2;R
RRRRRRRRR#PkLN5DRPkNDCN'sM2oCRR:=PkNDCR;
RRRRRRRRR0sCkRsM0#F_0MsHok5#LDPN2R;
RRRRRCRRD
#CRRRRRRRRRCRs0MksR_0F#H0sM5oRsHC#x5CRPkNDCP,RNCDk'oEHE-,R4;22
RRRRRRRR8CMR;HV
RRRRCRRD
#CRRRRRRRR#8HMG=R:R
4;RRRRRRRRVRFsHMRHRDPNkEC'HRoE8MFI0PFRNCDk'IDFRFDFbR
RRRRRRRRRHHVRR-=R4ER0CRM
RRRRRRRRR#RR5M#H8RG2:'=R3
';RRRRRRRRRRRR#8HMGRRRRR:=#8HMGRR+4R;
RRRRRRRRR8CMR;HV
RRRRRRRR#RR5M#H8RG2:v=Re_pg0OF_E5Ns1_a7ztpmQPB5NCDk52H22R;
RRRRRRRRRM#H8RGRR=R:RM#H8+GRR
4;RRRRRRRRCRM8DbFF;R
RRRRRRCRs0MksR
#;RRRRRMRC8VRH;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0F#H0sM
o;
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:z h)1emp k7_VCHG8s2RCs0kMaR1)tQhR
H#RRRRO#FM00NMRCDMRRR:Q hatR ):5=R-peqzD 'F.I+2;/d
RRRRsPNHDNLCkR#LDPNRz:Rh1) m pe7V_kH8GCRN5PD'kCEEHoRI8FMR0F-;d2
RRRRsPNHDNLCbRDN:8RR71a_mzpt_QBea Bm5)RjFR0RM5DCR*d+qRep'z D2FIR2-4;R
RRNRPsLHND#CRD:PRR71a_mzpt_QBea Bm5)RPkNDCC'DMEo0-84RF0IMF2Rj;R
RLHCoMR
RRVRHRDPNkDC'C0MoERR<4ER0CRM
RRRRR0sCkRsMh;z1
RRRR#CDCR
RRRRRHPVRNCDk'oEHERR<jER0CRM
RRRRRHRRVNRPD5kCPkNDCH'EoRE2=ZR''ER0CRM
RRRRRRRRR0sCkRsM0FF_#H0sM5oRsHC#x5CR#GVHCP85NCDk2.,R,NRPD'kCD2FI2R;
RRRRRCRRD
#CRRRRRRRRRCRs0MksR_0FFs#0HRMo5#sCHRxC5DPNkRC,.P,RNCDk'IDF2
2;RRRRRRRRCRM8H
V;RRRRRDRC#RHVPkNDCF'DI=R>R0jRE
CMRRRRRRRRHQVR#R_X5DPNkPC5NCDk'IDF202RE
CMRRRRRRRRRkR#LDPNRR:=5EF0CRs#=P>RNCDk5DPNkDC'F2I2;R
RRRRRRRRR#PkLN5DRPkNDCN'sM2oCRR:=PkNDCR;
RRRRRRRRR0sCkRsM0FF_#H0sM#o5kNLPD
2;RRRRRRRRCCD#
RRRRRRRRsRRCs0kMFR0_0F#soHMRC5s#CHxRN5PD,kCRDPNkEC'H,oER2-d2R;
RRRRRCRRMH8RVR;
RRRRR#CDCR
RRRRRRDR#P=R:R_0F#PkDRN5PD2kC;R
RRRRRRVRHR_Q#XPR5NCDkRN5PD'kCD2FI2ER0CRM
RRRRRRRRRNDb8=R:R05FE#CsRR=>PkNDCPR5NCDk'IDF2
2;RRRRRRRRCCD#
RRRRRRRRDRRbRN8:5=RFC0Es=#R>jR''
2;RRRRRRRRCRM8H
V;RRRRRRRRskC0s0MRF#_F0MsHoD5#PD5#PH'Eo8ERF0IMFDR#PH'EoeE-q pz'oEHE
22RRRRRRRRRRR&"
3"RRRRRRRRRRR&0FF_#H0sM#o5D#P5DEP'H-oEezqp H'Eo4E-RI8FMR0Fj&2RRNDb8
2;RRRRRMRC8VRH;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FFs#0H;Mo
R
RVOkM0MHFR_0FEs#0HRMo5DPNk:CRR)zh p1me_ 7kGVHCR82skC0s1MRah)Qt#RH
RRRRMOF#M0N0MRDC:RRRaQh )t RR:=5q-ep'z D+FIdc2/;R
RRNRPsLHND#CRkNLPDRR:z h)1emp k7_VCHG8PR5NCDk'oEHEFR8IFM0R2-c;R
RRNRPsLHNDDCRbRN8:aR17p_zmBtQ_Be aRm)50jRFDR5McC*Re+Rq pz'IDF24R-2R;
RPRRNNsHLRDC#RDP:aR17p_zmBtQ_Be aRm)5DPNkDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RHRRVNRPD'kCDoCM0<ERR04RE
CMRRRRRCRs0MksR1hz;R
RRDRC#RC
RRRRRRHVPkNDCH'Eo<ERR0jRE
CMRRRRRRRRHPVRNCDk5DPNkEC'H2oER'=RZ0'RE
CMRRRRRRRRRCRs0MksR_0FEs#0HRMo5#sCHRxC5H#VG5C8PkNDCR2,dP,RNCDk'IDF2
2;RRRRRRRRCCD#
RRRRRRRRsRRCs0kMFR0_0E#soHMRC5s#CHxRN5PD,kCRRd,PkNDCF'DI;22
RRRRRRRR8CMR;HV
RRRRCRRDV#HRDPNkDC'F>IR=RRj0MEC
RRRRRRRRRHVQX#_RN5PD5kCPkNDCF'DIR220MEC
RRRRRRRR#RRkNLPD=R:R05FE#CsRR=>PkNDCN5PD'kCD2FI2R;
RRRRRRRRRL#kPRND5DPNksC'NCMo2=R:RDPNk
C;RRRRRRRRRCRs0MksR_0FEs#0H5Mo#PkLN;D2
RRRRRRRR#CDCR
RRRRRRRRRskC0s0MRF#_E0MsHosR5Cx#HCPR5NCDk,NRPD'kCEEHo,cR-2
2;RRRRRRRRCRM8H
V;RRRRRDRC#RC
RRRRR#RRD:PR=FR0_D#kPPR5NCDk2R;
RRRRRHRRV#RQ_5XRPkNDCPR5NCDk'IDF202RE
CMRRRRRRRRRbRDN:8R=FR50sEC#>R=RDPNkPC5NCDk'IDF2
2;RRRRRRRRCCD#
RRRRRRRRDRRbRN8:5=RFC0Es=#R>jR''
2;RRRRRRRRCRM8H
V;RRRRRRRRskC0s0MRF#_E0MsHoD5#PD5#PH'Eo8ERF0IMFDR#PH'EoeE-q pz'oEHE
22RRRRRRRRRRR&"
3"RRRRRRRRRRR&0EF_#H0sM#o5D#P5DEP'H-oEezqp H'Eo4E-RI8FMR0FjD2&b2N8;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F0MRF#_E0MsHo
;
RkRVMHO0F0MRF#_F0MsHoPR5NCDkRz:Rh1) m pe7V_#H8GC2CRs0MksR)1aQRhtHR#
RORRF0M#NRM0MRCRRQ:Rhta  :)R=5R5PkNDCH'Eo4E+22+./
d;RRRRPHNsNCLDR8bNRRR:1_a7ztpmQeB_ mBa)R5j05FRMdC*R5-RPkNDCH'Eo4E+2-2RR;42
RRRRMOF#M0N0MRDC:RRRaQh )t RR:=5q-ep'z D+FI.d2/;R
RRNRPsLHND#CRkNLPDRR:z h)1emp #7_VCHG8PR5NCDk'oEHEFR8IFM0R2-d;R
RRNRPsLHNDDCRbRN8:aR17p_zmBtQ_Be aRm)50jRFDR5MdC*Re+Rq pz'IDF24R-2R;
RPRRNNsHLRDC#RDPR1:Raz7_pQmtB _eB)amRq5ep'z EEHoRe-Rq pz'IDFRI8FMR0Fj
2;RCRLo
HMRRRRHPVRNCDk'MDCoR0E<RR40MEC
RRRRsRRCs0kMzRh1R;
RCRRD
#CRRRRRVRHRDPNkEC'HRoE<RRj0MEC
RRRRRRRR0sCkRsM0FF_#H0sM5oRsHC#x5CRPkNDC.,R,NRPD'kCD2FI2R;
RRRRR#CDHPVRNCDk'IDFRR>=jER0CRM
RRRRRHRRV#RQ_5XRPkNDCN5PD'kCD2FI2ER0CRM
RRRRRRRRRL#kPRND:5=RFC0Es=#R>NRPD5kCPkNDCF'DI;22
RRRRRRRR#RRkNLPDPR5NCDk'MsNoRC2:P=RNCDk;R
RRRRRRRRRskC0s0MRF#_F0MsHok5#LDPN2R;
RRRRRCRRD
#CRRRRRRRRRCRs0MksR_0FFs#0HRMo5#sCHRxC5DPNkRC,PkNDCH'EoRE,-2d2;R
RRRRRRMRC8VRH;R
RRRRRCCD#
RRRRRRRR8bNRR:=5EF0CRs#=P>RNCDk5DPNkEC'H2oE2R;
RRRRR#RRD:PR=FR0_D#kPPR5NCDk2R;
RRRRRHRRV#RQ_5XRPkNDCPR5NCDk'IDF202RE
CMRRRRRRRRRbRDN:8R=FR50sEC#>R=RDPNkPC5NCDk'IDF2
2;RRRRRRRRCCD#
RRRRRRRRDRRbRN8:5=RFC0Es=#R>jR''
2;RRRRRRRRCRM8H
V;RRRRRRRRskC0s0MRF#_F0MsHoN5b8RR&#5DP#'DPEEHoRI8FMR0F#'DPEEHo-peqzE 'H2oE2R
RRRRRRRRR&3R""R
RRRRRRRRR&FR0_0F#soHM5P#D5P#D'oEHEq-ep'z EEHo-84RF0IMF2RjRD&Rb2N8;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F0MRF#_F0MsHo
;
RkRVMHO0F0MRF#_E0MsHoPR5NCDkRz:Rh1) m pe7V_#H8GC2CRs0MksR)1aQRhtHR#
RORRF0M#NRM0MRCRRQ:Rhta  :)R=5R5PkNDCH'Eo4E+22+d/
c;RRRRPHNsNCLDR8bNRRR:1_a7ztpmQeB_ mBa)R5j05FRMcC*R5-RPkNDCH'Eo4E+2-2RR;42
RRRRMOF#M0N0MRDC:RRRaQh )t RR:=5q-ep'z D+FIdc2/;R
RRNRPsLHND#CRkNLPDRR:z h)1emp #7_VCHG8PR5NCDk'oEHEFR8IFM0R2-c;R
RRNRPsLHNDDCRbRN8:aR17p_zmBtQ_Be aRm)50jRFDR5McC*Re+Rq pz'IDF24R-2R;
RPRRNNsHLRDC#RDPR1:Raz7_pQmtB _eB)amRN5PD'kCDoCM04E-RI8FMR0Fj
2;RCRLo
HMRRRRHPVRNCDk'MDCoR0E<RR40MEC
RRRRsRRCs0kMzRh1R;
RCRRD
#CRRRRRVRHRDPNkEC'HRoE<RRj0MEC
RRRRRRRR0sCkRsM0EF_#H0sM5oRsHC#x5CRPkNDCd,R,NRPD'kCD2FI2R;
RRRRR#CDHPVRNCDk'IDFRR>=jER0CRM
RRRRRHRRV#RQ_5XRPkNDCN5PD'kCD2FI2ER0CRM
RRRRRRRRRL#kPRND:5=RFC0Es=#R>NRPD5kCPkNDCF'DI;22
RRRRRRRR#RRkNLPDPR5NCDk'MsNoRC2:P=RNCDk;R
RRRRRRRRRskC0s0MRF#_E0MsHok5#LDPN2R;
RRRRRCRRD
#CRRRRRRRRRCRs0MksR_0FEs#0HRMo5#sCHRxC5DPNkRC,PkNDCH'EoRE,-2c2;R
RRRRRRMRC8VRH;R
RRRRRCCD#
RRRRRRRRP#DRR:=0#F_kRDP5DPNk;C2
RRRRRRRR8bNRR:=5EF0CRs#=P>RNCDk5DPNkEC'H2oE2R;
RRRRRHRRV#RQ_5XRPkNDCPR5NCDk'IDF202RE
CMRRRRRRRRRbRDN:8R=FR50sEC#>R=RDPNkPC5NCDk'IDF2
2;RRRRRRRRCCD#
RRRRRRRRDRRbRN8:5=RFC0Es=#R>jR''
2;RRRRRRRRCRM8H
V;RRRRRRRRskC0s0MRF#_E0MsHoN5b8RR&#5DP#'DPEEHoRI8FMR0F#'DPEEHo-peqzE 'H2oE2R
RRRRRRRRR&3R""R
RRRRRRRRR&FR0_0E#soHM5P#D5P#D'oEHEq-ep'z EEHo-84RF0IMF2RjRD&Rb2N8;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F0MRF#_E0MsHo
;
R-R-RFwsl0R#soHMRMVkOF0HMN#RDIDFRk$FRR0FOPFMCRs0N0R#soHMR0HMFRRNVCHG8R
R-b-RF0HMRlMkL3CsRGR NDlbCR:
RR--Ro#HMRNDkRV4:VRkH8GCRR5d8MFI0-FRd
2;R-R-RVRk4=R<RFVsl0_#soHMRj5"434j4"jj,VRk4H'EoRE,k'V4D2FI;-R-R6n3
-RR-ERaC3R""#RHR0FbHNFMDMRHRH0E#$R#MG0N,FREICCPs0RHRHCG#N0RMH8R#R
R-H-RMER0CsRIFRMoDNFO0MHFRRNMCFsss#RHRFbs8CkO8R3RmsPCVIDFRDIHDR
R-s-RCD#k0MRHR0#Nk0sNH3FM
VRRk0MOHRFMVlsF_s#0HRMo5R
RR#RL0MsHoRRRRRRRRRRRR:RRR)1aQ;htRRRRR-R-RMLHNRs$#H0sMRo
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)R;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDpCRRRRRRRR:p Qh;R
RRNRPsLHNDoCRFRF8RRR:Apmm ;qh
LRRCMoH
RRRR:pR=CRMIaR1)tQh'#5L0MsHo
2;RRRRs8CNR,5pR#sCk,D0RFoF8
2;RRRR8DCNDNFO05CRp
2;RRRRNC##s50Ro8FF2R
RRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR"&RVlsF_s#0H:MoR8ANRs#0HRMo"L&R#H0sM#oRCsPCHR0$CFsssR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRFVsl0_#soHM;R

RR--mNO0DMRN8CREGFROMsPC#MHF#FRIsN	R#FRVDIDF#R:
RR--kRV4<V=Rs_FlEs#0HRMo53"nUR",d-,RdR2;-n-R356RL0F0FxlRC#sFRF8sb8bC2R
R-k-RV<4R=sRVFFl_#H0sM5oR"3jncR",d-,RdR2;-n-R356R0RFbxFCs#sR8FCbb8R2
RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRRRRRRRRRRRRRR:1Qa)hRt;RRRRRR--mNO0D0R#soHM
RRRRMOF#M0N0CRDVH0_MG8CRRR:Q hat; )
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hat2 )
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7kGVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRRpRRRRR:QRph
 ;RRRRPHNsNCLDRFoF8RRR:mRAmqp hR;
RoLCHRM
RpRRRR:=MRCI1Qa)h5t'Fs#0H2Mo;R
RRsRFCRN85Rp,skC#DR0,o8FF2R;
R8RRCDNDF0ONCpR52R;
RNRR#s#C0oR5F2F8
RRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRR&VR"s_FlFs#0H:MoR8ANRs#0HRMo"F&R#H0sM#oRCsPCHR0$CFsssR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRFVsl#_F0MsHo
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHoRRRRRRRRRRRR:RRR)1aQ;htRRRRR-R-RGECRs#0H
MoRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp k7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCpRRRR:RRRhpQ R;
RPRRNNsHLRDCo8FFR:RRRmAmph q;R
RLHCoMR
RRRRp:M=RC1IRah)QtE'5#H0sM;o2
RRRRCEsN58Rps,RCD#k0o,RF2F8;R
RRCR8NFDDOCN0R25p;R
RR#RN#0CsRF5oF
82RRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRR&RRRs"VFEl_#H0sMRo:ARN8#H0sM"oR&#RE0MsHoCR#PHCs0C$RsssF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMVlsF_0E#soHM;R
R
VRRk0MOHRFMVlsF_s#0HRMo5R
RR#RL0MsHoRRRRRRRRRRRR:RRR)1aQ;htRRRRR-R-RMLHNRs$#H0sMRo
RORRF0M#NRM0D0CV_8HMCRGR:hRQa  t)R;
RORRF0M#NRM0sEHo0M_H8RCG:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _H#VG
C8R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7V_#H8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H82CG;R
RRNRPsLHNDpCRRRRRRRR:p Qh;R
RRNRPsLHNDoCRFRF8RRR:Apmm ;qh
LRRCMoH
RRRR:pR=CRMIaR1)tQh'#5L0MsHo
2;RRRRs8CNR,5pR#sCk,D0RFoF8
2;RRRR8DCNDNFO05CRp
2;RRRRNC##s50Ro8FF2R
RRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRR"&RVlsF_s#0H:MoR8ANRs#0HRMo"L&R#H0sM#oRCsPCHR0$CFsssR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRFVsl0_#soHM;R

RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRRRRRRRRRRRRRR:1Qa)hRt;RRRRRR--mNO0D0R#soHM
RRRRMOF#M0N0CRDVH0_MG8CRRR:Q hat; )
RRRRMOF#M0N0HRso_E0HCM8GRR:Q hat2 )
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8G
2;RRRRPHNsNCLDRRpRRRRR:QRph
 ;RRRRPHNsNCLDRFoF8RRR:mRAmqp hR;
RoLCHRM
RpRRRR:=MRCI1Qa)h5t'Fs#0H2Mo;R
RRsRFCRN85Rp,skC#DR0,o8FF2R;
R8RRCDNDF0ONCpR52R;
RNRR#s#C0oR5F2F8
RRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRR&VR"s_FlFs#0H:MoR8ANRs#0HRMo"F&R#H0sM#oRCsPCHR0$CFsssR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRFVsl#_F0MsHo
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHoRRRRRRRRRRRR:RRR)1aQ;htRRRRR-R-RGECRs#0H
MoRRRRO#FM00NMRVDC0M_H8RCGRQ:Rhta  
);RRRRO#FM00NMRosHEH0_MG8CRQ:Rhta  
)2RRRRskC0szMRh1) m pe7V_#H8GC
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp #7_VCHG8DR5C_V0HCM8GFR8IFM0RosHEH0_MG8C2R;
RPRRNNsHLRDCpRRRR:RRRhpQ R;
RPRRNNsHLRDCo8FFR:RRRmAmph q;R
RLHCoMR
RRRRp:M=RC1IRah)QtE'5#H0sM;o2
RRRRCEsN58Rps,RCD#k0o,RF2F8;R
RRCR8NFDDOCN0R25p;R
RR#RN#0CsRF5oF
82RRRRRCRsb0FsRGVHCb8_	Ho'MN#0M_OCMCNl
RRRR&RRRs"VFEl_#H0sMRo:ARN8#H0sM"oR&#RE0MsHoCR#PHCs0C$RsssF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMVlsF_0E#soHM;R

RR--1CNlRRN#NPLFC",R#CHx_#sC"#RHRCk#8FRVs0RH's#RNCMoRDFM$R3
VOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoR:aR1)tQh;RRRRRRRRRRRRRRRR-RR-HRLM$NsRs#0H
MoRRRR#CHx_#sCRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRFVsl0_#soHMR#5L0MsHo#,RH_xCs'C#EEHo,HR#xsC_CD#'F;I2
CRRMV8Rk0MOHRFMVlsF_s#0H;Mo
R
RVOkM0MHFRFVsl#_F0MsHo
R5RRRRFs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-m-ROD0NRs#0H
MoRRRR#CHx_#sCRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRFVsl#_F0MsHoFR5#H0sMRo,#CHx_#sC'oEHE#,RH_xCs'C#D2FI;R
RCRM8VOkM0MHFRFVsl#_F0MsHo
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHo:RRR)1aQ;htRRRRRRRRRRRRRRRRR-R-RGECRs#0H
MoRRRR#CHx_#sCRz:Rh1) m pe7V_kH8GC2R
RRCRs0MksR)zh p1me_ 7kGVHCH8R#R
RLHCoMR
RRCRs0MksRFVsl#_E0MsHo#5E0MsHo#,RH_xCs'C#EEHo,HR#xsC_CD#'F;I2
CRRMV8Rk0MOHRFMVlsF_0E#soHM;R

RMVkOF0HMsRVF#l_0MsHo
R5RRRRLs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-L-RHsMN$0R#soHM
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMsRVF#l_0MsHoLR5#H0sMRo,#CHx_#sC'oEHE#,RH_xCs'C#D2FI;R
RCRM8VOkM0MHFRFVsl0_#soHM;R

RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRR:1Qa)hRt;RRRRRRRRRRRRRRRRRR--mNO0D0R#soHM
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMsRVFFl_#H0sM5oRFs#0H,MoRx#HCC_s#H'EoRE,#CHx_#sC'IDF2R;
R8CMRMVkOF0HMsRVFFl_#H0sM
o;
VRRk0MOHRFMVlsF_0E#soHMRR5
RERR#H0sMRoR:aR1)tQh;RRRRRRRRRRRRRRRR-RR-CREG0R#soHM
RRRRx#HCC_s#RR:z h)1emp #7_VCHG8R2
RsRRCs0kMhRz)m 1p7e _H#VGRC8HR#
RoLCHRM
RsRRCs0kMsRVFEl_#H0sM5oREs#0H,MoRx#HCC_s#H'EoRE,#CHx_#sC'IDF2R;
R8CMRMVkOF0HMsRVFEl_#H0sM
o;
-RR-HR7s0CORMOFP#CsHRFMVOkM0MHF#R3R lGNb:DC
-RR-#RRHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-R-RkRV4<V=Rs_Fl#H0sM5oR"4j4jj34j;"2RR--n
36R-R-RRQM0#EHR#ONCER0C3R""#RHR0MFR0FbHNFMDN,RM08RE#CRHRxCFRV
RR--0RECFbk0kl0RkR#0lON0EGRCNDO0$R3
RR--bbksF:#CRDBNONkD00CRE#CR0MsHoFRLkNM8s#HC
bRRsCFO8CksRDONONkD0#C_0MsHoF_LksM8$
R5RRRRNRsoRRRRRRRR:MRHRaR1)tQh;RRRRRRRRRRR-H-RM0bkRs#0H
MoRRRRD0CV_8HMCRGR:kRF0hRQa  t)R;RRRRRRRRR-D-RC
V0RRRRsEHo0M_H8RCG:kRF0hRQa  t)H2R#RRRRRRR-s-RH0oE
RRRRR--ClGNb#DCRj"4j3j44"44RkIFDs8RCs0kMcR+,dR-
RRRRR--"Xj(3"ccRkIFDs8RCs0kM.R+,.R-RE50C0MREFCROD0NRksF0CHMRkIFDl8RkHD0b2D$
RRRRR--"Aq__B3_"FRIkRD8skC0s+MR4-,R40R5ERCM0RECERCGs0FkHRMCIDFk8kRlDb0HD
$2RRRRNNDH#NRGs:oRR)1aQRht5oNs'MDCoR0E8MFI04FR2#RHRoNs;-RR-NRl	HCR0FR8IFM0RMsNoRC
RPRRNNsHLRDCDs,RRQ:Rhta  R);RRRRRRRRR-RR-MRH0MCsNHDRMG8CCR#
RPRRNNsHLRDCVMFk808FRA:Rm mpq:hR=NRVD;#C
LRRCMoH
RRRRRHVN'soDoCM0>ERR0jRE
CMRRRRRRRD:G=RN'soEEHoR4-R;R
RRRRRs=R:R
j;RRRRRFRVsRRHHGMRN'sosoNMCFRDFRb
RRRRRHRRVNRGsHo52RR='R_'0MEC
RRRRRRRRHRRVRRs=RRj0MEC
RRRRRRRRRRRR:DR=RRD-;R4
RRRRRRRRCRRD
#CRRRRRRRRRRRRs=R:R+sRR
4;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVGoNs5RH2=RR''sRFRsGNo25HRh=RAR1uFGsRN5soH=2RRR]a0MEC
RRRRRRRRsRRCsbF0HRVG_C8b'	oH0M#NCMO_lMNCR
RRRRRRRRRRRR&"kwFMN8RRN#bOHCRMER0CMRHbRk01Qa)h"tRRG&RN
soRRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRCHD#VNRGsHo52RR='R3'0MEC
RRRRRRRRHRRVFRVk8M8F00RE
CMRRRRRRRRRRRRsFCbsV0RH8GC_ob	'#HM0ONMCN_MlRC
RRRRRRRRRRRRR"&RwMFk8IR0FHRLM$NsRHbFMR0#HHMRM0bkRs#0HRMo"RR&GoNs
RRRRRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR#CDCR
RRRRRRRRRRRRD:D=RRH-R;R
RRRRRRRRRRRRs:-=RHRR+4R;
RRRRRRRRRVRRF8kM8RF0:0=Rs;kC
RRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRVDC0M_H8RCG:D=R;R
RRRRRsEHo0M_H8RCG:s=R;R
RRDRC#RC
RRRRRVDC0M_H8RCG:j=R;R
RRRRRsEHo0M_H8RCG:j=R;R
RRMRC8VRH;R
RCRM8bOsFCs8kCNRODDOkN_0C#H0sMLo_F8kMs
$;
-RR-HR7s0CORMOFP#CsHRFMVOkM0MHF#R3R lGNb:DC
-RR-#RRHNoMDVRk4RR:kGVHC58RdFR8IFM0R2-d;R
R-R-RkRV4<V=Rs_Fl#H0sM5oR"4j4jj34j;"2RR--n
36R-R-RRQM0#EHR#ONCER0C3R""#RHR0MFR0FbHNFMDN,RM08RE#CRHRxCFRV
RR--0RECFbk0kl0RkR#0lON0EGRCNDO0$R3
RMVkOF0HMsRVF#l_0MsHo
R5RRRRLs#0HRMo:aR1)tQh2RRRRRRRRRRRRRRRRRRRR-RR-HRLM$NsRs#0H
MoRRRRskC0szMRh1) m pe7V_kH8GC
HRR#R
RRNRPsLHNDDCRC_V0HCM8Gs,RH0oE_8HMC:GRRaQh )t ;R
RLHCoMR
RRNRODDOkN_0C#H0sMLo_F8kMs5$RLs#0H,MoRVDC0M_H8,CGRosHEH0_MG8C2R;
RsRRCs0kMsRVF#l_0MsHoLR5#H0sMRo,D0CV_8HMCRG,sEHo0M_H82CG;R
RCRM8VOkM0MHFRFVsl0_#soHM;R

RR--7CHsOF0ROD0NR8NMRGECRMOFP#CsHRFMVOkM0MHF#R3RQ0MRERH#OCN#
-RR-ER0C0R#soHMRMDCo#0ER#lk0NRl03OERGR NDlbCR:
RR--#MHoN#DRV:4R=VR#H8GCRR568MFI0-FRd
2;R-R-R4#VRR<=VlsF_0F#soHMR(5"4"3c2-R-R3-n6R
RVOkM0MHFRFVsl#_F0MsHo
R5RRRRFs#0HRMo:aR1)tQh2RRRRRRRRRRRRRRRRRRRR-RR-ORm0RND#H0sMRo
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRsPNHDNLCCRDVH0_MG8C,HRso_E0HCM8GRR:Q hat; )
LRRCMoH
RRRRDONONkD0#C_0MsHoF_LksM8$FR5#H0sMRo,D0CV_8HMCRG,sEHo0M_H82CG;R
RRCRs0MksRFVsl#_F0MsHoFR5#H0sMRo,5C5DVH0_MG8C+*42d42-,HRso_E0HCM8G2*d;R
RCRM8VOkM0MHFRFVsl#_F0MsHo
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHoRR:1Qa)hRt2RRRRRRRRRRRRRRRRRRRRRR--ERCG#H0sMRo
RsRRCs0kMhRz)m 1p7e _HkVG
C8R#RH
RRRRsPNHDNLCCRDVH0_MG8C,HRso_E0HCM8GRR:Q hat; )
LRRCMoH
RRRRDONONkD0#C_0MsHoF_LksM8$ER5#H0sMRo,D0CV_8HMCRG,sEHo0M_H82CG;R
RRCRs0MksRFVsl#_E0MsHoER5#H0sMRo,5C5DVH0_MG8C+*42c42-,HRso_E0HCM8G2*c;R
RCRM8VOkM0MHFRFVsl#_E0MsHo
;
RkRVMHO0FVMRs_Fl#H0sM5oR
RRRR0L#soHMR1:Rah)QtR2RRRRRRRRRRRRRRRRRRRRR-L-RHsMN$0R#soHM
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCD0CV_8HMCRG,sEHo0M_H8RCG:hRQa  t)R;
RoLCHRM
RORRNkDODCN0_s#0H_MoLMFk8Rs$50L#soHM,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRskC0sVMRs_Fl#H0sM5oRLs#0H,MoRVDC0M_H8,CGRosHEH0_MG8C2R;
R8CMRMVkOF0HMsRVF#l_0MsHo
;
RkRVMHO0FVMRs_FlFs#0HRMo5R
RR#RF0MsHoRR:1Qa)hRt2RRRRRRRRRRRRRRRRRRRRRR--mNO0D0R#soHM
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCD0CV_8HMCRG,sEHo0M_H8RCG:hRQa  t)R;
RoLCHRM
RORRNkDODCN0_s#0H_MoLMFk8Rs$50F#soHM,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRskC0sVMRs_FlFs#0HRMo50F#soHM,5R5D0CV_8HMC4G+22*d-R4,sEHo0M_H8*CGd
2;RMRC8kRVMHO0FVMRs_FlFs#0H;Mo
R
RVOkM0MHFRFVsl#_E0MsHo
R5RRRREs#0HRMo:aR1)tQh2RRRRRRRRRRRRRRRRRRRR-RR-CREG0R#soHM
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCD0CV_8HMCRG,sEHo0M_H8RCG:hRQa  t)R;
RoLCHRM
RORRNkDODCN0_s#0H_MoLMFk8Rs$50E#soHM,CRDVH0_MG8C,HRso_E0HCM8G
2;RRRRskC0sVMRs_FlEs#0HRMo50E#soHM,5R5D0CV_8HMC4G+22*c-R4,sEHo0M_H8*CGc
2;RMRC8kRVMHO0FVMRs_FlEs#0H;Mo

RRR-R-RDs0_M#$0#ECHF#RMR
R-b-RslNoN$R#MC0E#_H#F
M
CRM8b	NONRoCL$F8RGVHCo8_CsMCHbO_	
o;
