7'h00: rv_rd_data = 32'h0080006f;
7'h01: rv_rd_data = 32'h12802623;
7'h02: rv_rd_data = 32'h7b349073;
7'h03: rv_rd_data = 32'h12002483;
7'h04: rv_rd_data = 32'h00905463;
7'h05: rv_rd_data = 32'h7b241073;
7'h06: rv_rd_data = 32'hf1402473;
7'h07: rv_rd_data = 32'h12802223;
7'h08: rv_rd_data = 32'h02848263;
7'h09: rv_rd_data = 32'h4004c493;
7'h0a: rv_rd_data = 32'h00848663;
7'h0b: rv_rd_data = 32'h12002483;
7'h0c: rv_rd_data = 32'hff1ff06f;
7'h0d: rv_rd_data = 32'h12802423;
7'h0e: rv_rd_data = 32'h7b202473;
7'h0f: rv_rd_data = 32'h7b3024f3;
7'h10: rv_rd_data = 32'h7b200073;
7'h11: rv_rd_data = 32'h12902023;
7'h12: rv_rd_data = 32'h7b202473;
7'h13: rv_rd_data = 32'h7b3024f3;
7'h14: rv_rd_data = 32'h10000067;
