--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb/oIlbNbC/s#GHHDMDG/HoL/CsMCHoO/CoM_CsMCHsO/Nsl_IPb3E48yR-f
--

--
-
R--1bHlD)CRqIvRHR0E#oHMDqCR7 7)1V1RFLsRFR0Es8CNR8NMRHIs0-C
-NRas0oCRX:RHMDHG-
-
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;CHM00)$Rq)v_WHuR#o
SCsMCH5OR
VSSNDlH$RR:#H0sM:oR=MR"F"MC;S
SI0H8ERR:HCM0oRCs:.=R;SR
S8N8s8IH0:ERR0HMCsoCRR:=UR;RRRRRR-R-RoLHRFCMkRoEVRFs80CbES
S80CbERR:HCM0oRCs:.=R6
n;SFS8ks0_C:oRRFLFDMCNRR:=V#NDCR;RR-RR-NRE#kRF00bkRosC
8SSHsM_C:oRRFLFDMCNRR:=V#NDCR;RRRRR-E-RN8#RNR0NHkMb0CRsoS
SNs88_osCRL:RFCFDN:MR=NRVDR#CRRRRRR--ERN8Ns88CR##s
CoS;S2
FSbs50R
7SSm:zaR0FkR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
7SSQRhR:MRHR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2
qSS7R7):MRHR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2
WSS :RRRRHM#_08DHFoOR;RRRRRRR--I0sHCMRCNCLDRsVFRlsN
BSSp:iRRRHM#_08DHFoOR;RRRRRRR--OODF	FRVsNRslN,R8,8sRM8H
mSSBRpi:MRHR8#0_oDFHRORRRRRRR--FRb0OODF	FRVsFR8kS0
S
2;CRM8CHM00)$Rq)v_W
u;

---w-RH0s#RbHlDCClM00NHRFMl0k#RRLCODNDCN8RsjOE

--NEsOHO0C0CksRFLDOs	_NFlRVqR)vW_)u#RH
b0$CMRH0s_NsRN$HN#Rs$sNRR5j06FR2VRFR0HMCsoC;F
OMN#0MI0RHE80_sNsN:$RR0HM_sNsN:$R=4R5,,R.RRc,g4,RUd,Rn
2;O#FM00NMRb8C0NE_s$sNRH:RMN0_s$sNRR:=5d4nURc,U.4g,jRcgRn,.Ujc,jR4.Rc,624.;F
OMN#0M80RH.PdRH:RMo0CC:sR=IR5HE80-/42d
n;O#FM00NMRP8H4:nRR0HMCsoCRR:=58IH04E-2U/4;F
OMN#0M80RHRPU:MRH0CCos=R:RH5I8-0E4g2/;F
OMN#0M80RHRPc:MRH0CCos=R:RH5I8-0E4c2/;F
OMN#0M80RHRP.:MRH0CCos=R:RH5I8-0E4.2/;F
OMN#0M80RHRP4:MRH0CCos=R:RH5I8-0E442/;O

F0M#NRM0LDFF4RR:LDFFCRNM:5=R84HPRj>R2O;
F0M#NRM0LDFF.RR:LDFFCRNM:5=R8.HPRj>R2O;
F0M#NRM0LDFFcRR:LDFFCRNM:5=R8cHPRj>R2O;
F0M#NRM0LDFFURR:LDFFCRNM:5=R8UHPRj>R2O;
F0M#NRM0LDFF4:nRRFLFDMCNRR:=5P8H4>nRR;j2
MOF#M0N0FRLF.DdRL:RFCFDN:MR=8R5H.PdRj>R2
;
O#FM00NMRP8H4UndcRR:HCM0oRCs:5=R80CbE2-4/d4nU
c;O#FM00NMRP8HU.4gRH:RMo0CC:sR=8R5CEb0-/42U.4g;F
OMN#0M80RHjPcg:nRR0HMCsoCRR:=5b8C04E-2j/cg
n;O#FM00NMRP8H.UjcRH:RMo0CC:sR=8R5CEb0-/42.Ujc;F
OMN#0M80RHjP4.:cRR0HMCsoCRR:=5b8C04E-2j/4.
c;O#FM00NMRP8H6R4.:MRH0CCos=R:RC58b-0E462/4
.;
MOF#M0N0FRLF4D6.RR:LDFFCRNM:5=R86HP4>.RR;j2
MOF#M0N0FRLFjD4.:cRRFLFDMCNRR:=5P8H4cj.Rj>R2O;
F0M#NRM0LDFF.UjcRL:RFCFDN:MR=8R5HjP.c>URR;j2
MOF#M0N0FRLFjDcg:nRRFLFDMCNRR:=5P8HcnjgRj>R2O;
F0M#NRM0LDFFU.4gRL:RFCFDN:MR=8R5H4PUg>.RR;j2
MOF#M0N0FRLFnD4dRUc:FRLFNDCM=R:RH58Pd4nU>cRR;j2
F
OMN#0M#0RkIl_HE80RH:RMo0CC:sR=mRAmqp hF'b#F5LF2D4RA+Rm mpqbh'FL#5F.FD2RR+Apmm 'qhb5F#LDFFc+2RRmAmph q'#bF5FLFDRU2+mRAmqp hF'b#F5LFnD42O;
F0M#NRM0#_kl80CbERR:HCM0oRCs:6=RR5-RApmm 'qhb5F#LDFF624.RA+Rm mpqbh'FL#5F4FDj2.cRA+Rm mpqbh'FL#5F.FDj2cURA+Rm mpqbh'FL#5FcFDj2gnRA+Rm mpqbh'FL#5FUFD42g.2
;
O#FM00NMROI_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_RIOHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lH_I820E;F
OMN#0M80R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5k8l_CEb02O;
F0M#NRM08E_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_kl80CbE
2;
MOF#M0N0_RII0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E4I2/_FOEH_OCI0H8ERR+4O;
F0M#NRM0IC_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/OI_EOFHCC_8bR0E+;R4
F
OMN#0M80R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/428E_OFCHO_8IH0+ERR
4;O#FM00NMR88_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/8OHEFO8C_CEb0R4+R;O

F0M#NRM0IH_#x:CRR0HMCsoCRR:=IH_I8_0EM_klODCD#RR*IC_8b_0EM_klODCD#O;
F0M#NRM08H_#x:CRR0HMCsoCRR:=8H_I8_0EM_klODCD#RR*8C_8b_0EM_klODCD#
;
O#FM00NMRFLFDR_8:FRLFNDCM=R:R_58#CHxRI-R_x#HC=R<R;j2
MOF#M0N0FRLFID_RL:RFCFDN:MR=FRM0F5LF8D_2
;
O#FM00NMRFOEH_OCI0H8ERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OCI0H8E
2;O#FM00NMRFOEH_OC80CbERR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*_R8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IRI*R_FOEH_OC80CbE
2;O#FM00NMR8IH0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R58IH04E-2_/8OHEFOIC_HE802RR+5mAmph q'#bF5FLFD2_IR5*RI0H8E2-4/OI_EOFHCH_I820ER4+R;F
OMN#0M80RCEb0_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*5CEb0-/428E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RRC58b-0E4I2/_FOEH_OC80CbE+2RR
4;-F-OMN#0MM0RkOl_C#DDRH:RMo0CC:sR=5R55b8C0-ERRR42/.Rd2RR+5855CEb0R4-R2FRl8.Rd2RR/42n2;RRR-y-RRRFV)dqv.1X4RDOCDM#RCCC88-R
-MOF#M0N0CRDVF0_PRCs:MRH0CCos=R:R55580CbERR+4R62lRF8dR.2/nR42R;RRRRRRRRRRRRRRRRRRRRRR-RR-RRyF)VRqnv4XR41M8CCCV8RFDsRCRV0FsPCRsIF80#
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L.k#RF:RkL0_k_#.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#U0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjU,R*8IH0ME_kOl_C#DD+8(RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:URR0Fk_#LkU$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,.H*I8_0EM_klODCD#R+48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#R4n:NRbs$H0_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,dI.*HE80_lMk_DOCDd#+4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lkd:.RR0Fk_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_d.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lkd:.RRsbNH_0$Ldk#.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FINs88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRsN8C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RR--0sFRC#oH0RCs0REC#CCDO#0RHNoMDVRFRH0s#00NC0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjjjjjRj"&8RN_osC5;j2
MSC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjj"jjRN&R8C_soR548MFI0jFR2S;
CRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjjjjj"RR&Ns8_C.o5RI8FMR0Fj
2;S8CMRMoCC0sNC.Rz;R
RRdRzRRR:H5VRNs88I0H8ERR=co2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjj"RR&Ns8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjj"jjRN&R8C_soR5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80Rn=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjjjjj&"RR_N8s5Co6FR8IFM0R;j2
MSC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjRj"&8RN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFNI_8R8s<"=RjjjjjRj"&8RN_osC58(RF0IMF2Rj;C
SMo8RCsMCNR0Cz
(;RRRRzRUR:VRHR85N8HsI8R0E=2RgRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjj&"RR_N8s5CoUFR8IFM0R;j2
MSC8CRoMNCs0zCRUR;
RzRRg:RRRRHV58N8s8IH0=ERR24jRMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjj"RR&Ns8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFNI_8R8s<"=Rj"jjRN&R8C_soj54RI8FMR0Fj
2;S8CMRMoCC0sNC4RzjR;
RzRR4R4R:VRHR85N8HsI8R0E=.R42CRoMNCs0SC
RRRRD_FINs88RR<=""jjRN&R8C_so454RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz4R;
RzRR4R.R:VRHR85N8HsI8R0E=dR42CRoMNCs0SC
RRRRD_FINs88RR<='Rj'&8RN_osC5R4.8MFI0jFR2S;
CRM8oCCMsCN0R.z4;R
RR4Rzd:RRRRHV58N8s8IH0>ERR24dRMoCC0sNCR
SRDRRFNI_8R8s<N=R8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR-Q-RV8R5F_k0s2CoRosCHC#0smR7zkaR#oHMRpmBiR
RR4Rzn:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_CRo2LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRRzR4(RH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_soH5I8-0E4FR8IFM0R;j2
MSC8CRoMNCs0zCR4
(;
RRRRR--Q5VRNs88_osC2CRso0H#CqsR7R7)kM#HopRBi-
-RRRRzR4nRH:RVNR58_8ss2CoRMoCC0sNC-
-RRRRRRRRbOsFCR##5iBp,7Rq7R)2LHCoM-
-RRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EM-
-RRRRRRRRRRRRRRRRNs8_C<oR=7Rq7N)58I8sHE80-84RF0IMF2Rj;-
-RRRRRRRRRRRRCRM8H
V;-R-RRRRRRMRC8sRbF#OC#-;
-MSC8CRoMNCs0zCR4
n;-R-RR4Rz(RR:H5VRMRF0Ns88_osC2CRoMNCs0RC
RRRRRRRRRNRR8C_so=R<R7q7)-;
-MSC8CRoMNCs0zCR4
(;SRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1S4
zR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERRR4c2CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFcR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRc
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR4g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RcM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:jRRRHV58N8s8IH0>ERR24cRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjS;
-Q-RVNR58I8sHE80RR<=4Rc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.Rz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_d4nU4cXRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_d4nU4cXR):Rq4vAn4_1
RSRRRRRRRRRRFRbsl0RN5bR7jQ52>R=R_HMs5Co[R2,q)77RR=>D_FINs885R4d8MFI0jFR2 ,Rh>R=R''4,1R1)>R=R''j,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,7jm52>R=R0Fk_#Lk4,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_k5#4H2,[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;..
RRRRCRSMo8RCsMCNR0Cz;4g
RRRR8CMRMoCC0sNC4RzUR;RRRR
RRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1S.
zR.d:VRHRE5OFCHO_8IH0=ERRR.2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR24dRMoCC0sNCR
RRRRRRORzDR	:bOsFCR##5iBp2R
SRRRRRoLCHSM
RRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RSRRRRRRRRRNC8so85N8HsI8-0E4FR8IFM0R24dRR<=Ns8_CNo58I8sHE80-84RF0IMFdR42S;
SRRRCRM8H
V;SMSC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRS.:cRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>dR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.Sz6RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNC8so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0F4Rd2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6z.;-
S-VRQR85N8HsI8R0E<4=RdM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:nRRRHV58N8s8IH0<ER=dR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnz.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qvU.4gX:.RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAqUv_4Xg..RR:)Aqv41n_.R
SRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)>R=RIDF_8N8s.54RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4=2R>kRF0k_L#H.5,[.*+,42R57mj=2R>kRF0k_L#H.5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5[.*2=R<R0Fk_#Lk.,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5.[2+4RR<=F_k0L.k#5.H,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(z.;R
RRSRRCRM8oCCMsCN0Rcz.;R
RRMRC8CRoMNCs0zCR.Rd;RS

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHR85N8HsI8R0E>.R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF.R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR.
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.g:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R.M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:jRRRHV58N8s8IH0>ERR24.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24.RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRzjS;
-Q-RVNR58I8sHE80RR<=4R.2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRd4:VRHR85N8HsI8R0E<4=R.o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjnRXc:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvcnjgX:cRRv)qA_4n1Sc
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cco5*d[+RI8FMR0Fc2*[,7Rq7=)R>FRDI8_N84s54FR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75Rd2=F>RkL0_k5#cHc,R*d[+27,Rm25.RR=>F_k0Lck#5cH,*.[+2
,RSSSS74m52>R=R0Fk_#Lkc,5Hc+*[4R2,7jm52>R=R0Fk_#Lkc,5HR[c*2
2;RRRRRRRRRRRRRRRRF_k0s5Coc2*[RR<=F_k0Lck#5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R42<F=RkL0_k5#cH*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+.RR<=F_k0Lck#5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*d[+2=R<R0Fk_#Lkc,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1gSdzdRH:RVOR5EOFHCH_I8R0E=2RgRMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>4R42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMF4R42=R<R_N8s5CoNs88I0H8ER-48MFI04FR4
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R244RH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCdRz6S;
-Q-RVNR58I8sHE80RR<=4R42MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRdn:VRHR85N8HsI8R0E<4=R4o2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_c.jURXU:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv.UjcX:URRv)qA_4n1Sg
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_Cgo5*([+RI8FMR0Fg2*[,7Rq7=)R>FRDI8_N84s5jFR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R(2=F>RkL0_k5#UH*,U[2+(,mR75Rn2=F>RkL0_k5#UH*,U[2+n,SR
S7SSm256RR=>F_k0LUk#5UH,*6[+27,Rm25cRR=>F_k0LUk#5UH,*c[+27,Rm25dRR=>F_k0LUk#5UH,*d[+2
,RSSSS7.m52>R=R0Fk_#LkU,5HU+*[.R2,74m52>R=R0Fk_#LkU,5HU+*[4R2,7jm52>R=R0Fk_#LkU,5HU2*[,SR
S7SSQju52>R=R_HMs5Cog+*[UR2,75muj=2R>NRbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,2R[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;d(
RRRRCRSMo8RCsMCNR0Cz;dc
RRRR8CMRMoCC0sNCdRzd
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_4SU
zRdU:VRHRE5OFCHO_8IH0=ERR24URMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>jR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRj<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;j2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgzdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rj2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRcj:VRHR85N8HsI8R0E>jR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFjR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRc
j;SR--Q5VRNs88I0H8E=R<R24jRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zcRH:RVNR58I8sHE80RR<=4Rj2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRc
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSc:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_4.4cXnRR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_4.4cXnRR:)Aqv41n_4SU
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_C4o5U+*[486RF0IMFUR4*,[2R7q7)>R=RIDF_8N8sR5g8MFI0jFR2 ,Rh>R=R''4,1R1)>R=R''j,SR
SWSS >R=R0Is_5CMHR2,BRpi=B>RpRi,74m56=2R>kRF0k_L#54nHn,4*4[+6R2,74m5c=2R>kRF0k_L#54nHn,4*4[+cR2,
SSSS57m4Rd2=F>RkL0_kn#454H,n+*[4,d2R57m4R.2=F>RkL0_kn#454H,n+*[4,.2R57m4R42=F>RkL0_kn#454H,n+*[4,42RS
SSmS7524jRR=>F_k0L4k#n,5H4[n*+24j,mR75Rg2=F>RkL0_kn#454H,n+*[gR2,7Um52>R=R0Fk_#Lk4Hn5,*4n[2+U,S
SSmS75R(2=F>RkL0_kn#454H,n+*[(R2,7nm52>R=R0Fk_#Lk4Hn5,*4n[2+n,mR75R62=F>RkL0_kn#454H,n+*[6
2,SRSSR7RRm25cRR=>F_k0L4k#n,5H4[n*+,c2R57md=2R>kRF0k_L#54nHn,4*d[+27,Rm25.RR=>F_k0L4k#n,5H4[n*+,.2
RSSRRRRR7RRm254RR=>F_k0L4k#n,5H4[n*+,42R57mj=2R>kRF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_soU54*4[+(FR8IFM0R*4U[n+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5R42=b>RN0sH$k_L#54nH.,R*4[+27,Rmju52>R=RsbNH_0$L4k#n,5HR[.*2
2;RRRRRRRRRRRRRRRRF_k0s5Co4[U*2=R<R0Fk_#Lk4Hn5,*4n[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R42<F=RkL0_kn#454H,n+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R.2<F=RkL0_kn#454H,n+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rd2<F=RkL0_kn#454H,n+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rc2<F=RkL0_kn#454H,n+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R62<F=RkL0_kn#454H,n+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rn2<F=RkL0_kn#454H,n+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+R(2<F=RkL0_kn#454H,n+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+RU2<F=RkL0_kn#454H,n+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+Rg2<F=RkL0_kn#454H,n+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24jRR<=F_k0L4k#n,5H4[n*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+4<2R=kRF0k_L#54nHn,4*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24.RR<=F_k0L4k#n,5H4[n*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+d<2R=kRF0k_L#54nHn,4*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24cRR<=F_k0L4k#n,5H4[n*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+6<2R=kRF0k_L#54nHn,4*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24nRR<=bHNs0L$_kn#45.H,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[(+42=R<RsbNH_0$L4k#n,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCcRz.R;
RRRRS8CMRMoCC0sNCdRzgR;
RCRRMo8RCsMCNR0Cz;dU
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_n1d
cSzdRR:H5VROHEFOIC_HE80Rd=Rno2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVRR5Ns88I0H8ERR>gRR2oCCMsCN0
RSRRORzDR	:bOsFCR##5iBp2S
SRCRLo
HMSRSRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
SRRRRNRR8osC58N8s8IH04E-RI8FMR0Fg<2R=8RN_osC58N8s8IH04E-RI8FMR0Fg
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	S;
RRRRzRcc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzRc6:VRHR85N8HsI8R0E>2RgRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8S
SSkSF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECR85N_osC58N8s8IH04E-RI8FMR0Fg=2RRRH2CCD#R''j;S
SS8CMRMoCC0sNCcRz6S;
-Q-RVNR58I8sHE80RR<=gM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8SzSSc:nRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0Rnzc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSSc:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_6..XdRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRRRRRRRRRqA)v4_6..XdR):Rq4vAnd_1nR
RRRRRRRRRRRRRRRRRRFRbsl0RN5bR7=QR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7R7)=F>DI8_N8Us5RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRW =I>RsC0_M25H,pRBi>R=RiBp,mR752d4RR=>F_k0Ldk#.,5Hd[.*+2d4,mR752djRR=>F_k0Ldk#.,5Hd[.*+2dj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5g=2R>kRF0k_L#5d.H.,d*.[+gR2,7.m5U=2R>kRF0k_L#5d.H.,d*.[+UR2,7.m5(=2R>kRF0k_L#5d.H.,d*.[+(
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.nRR=>F_k0Ldk#.,5Hd[.*+2.n,mR752.6RR=>F_k0Ldk#.,5Hd[.*+2.6,mR752.cRR=>F_k0Ldk#.,5Hd[.*+2.c,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m5d=2R>kRF0k_L#5d.H.,d*.[+dR2,7.m5.=2R>kRF0k_L#5d.H.,d*.[+.R2,7.m54=2R>kRF0k_L#5d.H.,d*.[+4
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR752.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7524gRR=>F_k0Ldk#.,5Hd[.*+24g,mR7524URR=>F_k0Ldk#.,5Hd[.*+24U,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR74m5(=2R>kRF0k_L#5d.H.,d*4[+(R2,74m5n=2R>kRF0k_L#5d.H.,d*4[+nR2,74m56=2R>kRF0k_L#5d.H.,d*4[+6
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7524cRR=>F_k0Ldk#.,5Hd[.*+24c,mR7524dRR=>F_k0Ldk#.,5Hd[.*+24d,mR7524.RR=>F_k0Ldk#.,5Hd[.*+24.,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4R42=F>RkL0_k.#d5dH,.+*[4,42R57m4Rj2=F>RkL0_k.#d5dH,.+*[4,j2R57mg=2R>kRF0k_L#5d.H.,d*g[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75RU2=F>RkL0_k.#d5dH,.+*[UR2,7(m52>R=R0Fk_#LkdH.5,*d.[2+(,mR75Rn2=F>RkL0_k.#d5dH,.+*[nR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm256RR=>F_k0Ldk#.,5Hd[.*+,62R57mc=2R>kRF0k_L#5d.H.,d*c[+27,Rm25dRR=>F_k0Ldk#.,5Hd[.*+,d2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7.m52>R=R0Fk_#LkdH.5,*d.[2+.,mR75R42=F>RkL0_k.#d5dH,.+*[4R2,7jm52>R=R0Fk_#LkdH.5,*d.[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQ=uR>MRH_osC5*dn[6+dRI8FMR0Fd[n*+2d.,mR7u25dRR=>bHNs0L$_k.#d5RH,c+*[d
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u25.RR=>bHNs0L$_k.#d5RH,c+*[.R2,75mu4=2R>NRbs$H0_#LkdH.5,*Rc[2+4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75muj=2R>NRbs$H0_#LkdH.5,*Rc[;22
RRRRRRRRRRRRRRRRFRRks0_Cdo5n2*[RR<=F_k0Ldk#.,5Hd[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+4RR<=F_k0Ldk#.,5Hd[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.<2R=kRF0k_L#5d.H.,d*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+dRR<=F_k0Ldk#.,5Hd[.*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[c<2R=kRF0k_L#5d.H.,d*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+6RR<=F_k0Ldk#.,5Hd[.*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[n<2R=kRF0k_L#5d.H.,d*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+(RR<=F_k0Ldk#.,5Hd[.*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[U<2R=kRF0k_L#5d.H.,d*U[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[2+gRR<=F_k0Ldk#.,5Hd[.*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rj2<F=RkL0_k.#d5dH,.+*[4Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R42<F=RkL0_k.#d5dH,.+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R.2<F=RkL0_k.#d5dH,.+*[4R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rd2<F=RkL0_k.#d5dH,.+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rc2<F=RkL0_k.#d5dH,.+*[4Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R62<F=RkL0_k.#d5dH,.+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rn2<F=RkL0_k.#d5dH,.+*[4Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4R(2<F=RkL0_k.#d5dH,.+*[4R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4RU2<F=RkL0_k.#d5dH,.+*[4RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[4Rg2<F=RkL0_k.#d5dH,.+*[4Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rj2<F=RkL0_k.#d5dH,.+*[.Rj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R42<F=RkL0_k.#d5dH,.+*[.R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R.2<F=RkL0_k.#d5dH,.+*[.R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rd2<F=RkL0_k.#d5dH,.+*[.Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rc2<F=RkL0_k.#d5dH,.+*[.Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R62<F=RkL0_k.#d5dH,.+*[.R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rn2<F=RkL0_k.#d5dH,.+*[.Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.R(2<F=RkL0_k.#d5dH,.+*[.R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.RU2<F=RkL0_k.#d5dH,.+*[.RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[.Rg2<F=RkL0_k.#d5dH,.+*[.Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRj2<F=RkL0_k.#d5dH,.+*[dRj2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR42<F=RkL0_k.#d5dH,.+*[dR42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dR.2<b=RN0sH$k_L#5d.H*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*d[+d<2R=NRbs$H0_#LkdH.5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRc2<b=RN0sH$k_L#5d.H*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d6RR<=bHNs0L$_k.#d5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SMSC8CRoMNCs0zCRc
(;SMSC8CRoMNCs0zCRc
c;S8CMRMoCC0sNCcRzdC;
MN8RsHOE00COkRsCLODF	N_sl
;
-M-RFI_s_COEOV	RF#sRHDMoCFRbs)0RqHvR#8RHCHM0ORND0LFRD	FORlsN
ONsECH0Os0kCFRM__sIOOEC	VRFRv)q_u)WR
H#Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FMVRFI_s_COEO:	RRONsECH0Os0kC#RHR#"zHRMoLODF	N_slFRVsHR#MCoDRsbF0NRslHRI0#ER$sM_N0l#$RDCMsF_IE_OC"O	;$
0bHCRMN0_s$sNRRH#NNss$jR5RR0F6F2RVMRH0CCosO;
F0M#NRM0I0H8Es_NsRN$:MRH0s_NsRN$:5=R4.,R,,RcRRg,4RU,d;n2
MOF#M0N0CR8b_0ENNss$RR:H_M0NNss$=R:Rn54d,UcRgU4.c,Rj,gnRc.jU4,Rj,.cR.642O;
F0M#NRM08dHP.RR:HCM0oRCs:5=RI0H8E2-4/;dn
MOF#M0N0HR8PR4n:MRH0CCos=R:RH5I8-0E442/UO;
F0M#NRM08UHPRH:RMo0CC:sR=IR5HE80-/42gO;
F0M#NRM08cHPRH:RMo0CC:sR=IR5HE80-/42cO;
F0M#NRM08.HPRH:RMo0CC:sR=IR5HE80-/42.O;
F0M#NRM084HPRH:RMo0CC:sR=IR5HE80-/424
;
O#FM00NMRFLFD:4RRFLFDMCNRR:=5P8H4RR>j
2;O#FM00NMRFLFD:.RRFLFDMCNRR:=5P8H.RR>j
2;O#FM00NMRFLFD:cRRFLFDMCNRR:=5P8HcRR>j
2;O#FM00NMRFLFD:URRFLFDMCNRR:=5P8HURR>j
2;O#FM00NMRFLFDR4n:FRLFNDCM=R:RH58PR4n>2Rj;F
OMN#0ML0RFdFD.RR:LDFFCRNM:5=R8dHP.RR>j
2;
MOF#M0N0HR8Pd4nU:cRR0HMCsoCRR:=5b8C04E-2n/4d;Uc
MOF#M0N0HR8PgU4.RR:HCM0oRCs:5=R80CbE2-4/gU4.O;
F0M#NRM08cHPjRgn:MRH0CCos=R:RC58b-0E4c2/j;gn
MOF#M0N0HR8Pc.jURR:HCM0oRCs:5=R80CbE2-4/c.jUO;
F0M#NRM084HPjR.c:MRH0CCos=R:RC58b-0E442/j;.c
MOF#M0N0HR8P.64RH:RMo0CC:sR=8R5CEb0-/426;4.
F
OMN#0ML0RF6FD4:.RRFLFDMCNRR:=5P8H6R4.>2Rj;F
OMN#0ML0RF4FDjR.c:FRLFNDCM=R:RH58P.4jcRR>j
2;O#FM00NMRFLFDc.jURR:LDFFCRNM:5=R8.HPjRcU>2Rj;F
OMN#0ML0RFcFDjRgn:FRLFNDCM=R:RH58PgcjnRR>j
2;O#FM00NMRFLFDgU4.RR:LDFFCRNM:5=R8UHP4Rg.>2Rj;F
OMN#0ML0RF4FDncdURL:RFCFDN:MR=8R5HnP4dRUc>2Rj;O

F0M#NRM0#_klI0H8ERR:HCM0oRCs:A=Rm mpqbh'FL#5F4FD2RR+Apmm 'qhb5F#LDFF.+2RRmAmph q'#bF5FLFDRc2+mRAmqp hF'b#F5LF2DURA+Rm mpqbh'FL#5F4FDn
2;O#FM00NMRl#k_b8C0:ERR0HMCsoCRR:=6RR-5mAmph q'#bF5FLFD.642RR+Apmm 'qhb5F#LDFF4cj.2RR+Apmm 'qhb5F#LDFF.Ujc2RR+Apmm 'qhb5F#LDFFcnjg2RR+Apmm 'qhb5F#LDFFU.4g2
2;
MOF#M0N0_RIOHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lH_I820E;F
OMN#0MI0R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5kIl_HE802O;
F0M#NRM08E_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_kl80CbE
2;O#FM00NMRO8_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_b8C0;E2
F
OMN#0MI0R_8IH0ME_kOl_C#DDRH:RMo0CC:sR=IR5HE80-/42IE_OFCHO_8IH0+ERR
4;O#FM00NMR8I_CEb0_lMk_DOCD:#RR0HMCsoCRR:=5b8C04E-2_/IOHEFO8C_CEb0R4+R;O

F0M#NRM08H_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/O8_EOFHCH_I8R0E+;R4
MOF#M0N0_R880CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E482/_FOEH_OC80CbERR+4
;
O#FM00NMR#I_HRxC:MRH0CCos=R:RII_HE80_lMk_DOCD*#RR8I_CEb0_lMk_DOCD
#;O#FM00NMR#8_HRxC:MRH0CCos=R:RI8_HE80_lMk_DOCD*#RR88_CEb0_lMk_DOCD
#;
MOF#M0N0FRLF8D_RL:RFCFDN:MR=8R5_x#HCRR-IH_#x<CR=2Rj;F
OMN#0ML0RF_FDIRR:LDFFCRNM:M=RFL05F_FD8
2;
MOF#M0N0EROFCHO_8IH0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_8IH0;E2
MOF#M0N0EROFCHO_b8C0:ERR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8R8*R_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*IE_OFCHO_b8C0;E2
MOF#M0N0HRI8_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*H5I8-0E482/_FOEH_OCI0H8E+2RRm5Amqp hF'b#F5LFID_2RR*58IH04E-2_/IOHEFOIC_HE802RR+4O;
F0M#NRM080CbEk_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*80CbE2-4/O8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*8R5CEb0-/42IE_OFCHO_b8C0RE2+;R4
O--F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5C58bR0E-2R4Rd/R.+2RR55580CbERR-4l2RFd8R./2RR24n2R;RRR--yVRFRv)qd4.X1CRODRD#M8CCC
8R-F-OMN#0MD0RC_V0FsPCRH:RMo0CC:sR=5R55b8C0+ERR246R8lFR2d.R4/RnR2;RRRRRRRRRRRRRRRRRRRRRRRR-y-RRRFV)4qvn1X4RCMC8RC8VRFsD0CVRCFPsFRIs
8#0C$bR0Fk_#Lk4$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:4RR0Fk_#Lk4$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lkc$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0Lck#RF:RkL0_k_#c0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#0U_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,HRI8_0EM_klODCD#R-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#:URRsbNH_0$LUk#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,nR4*8IH0ME_kOl_C#DD+R468MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#4RF:RkL0_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRI.*HE80_lMk_DOCD4#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_kn#4Rb:RN0sH$k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFV80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Is_RCM:0R#8F_Do_HOP0COF8s5CEb0_lMk_DOCD4#-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDMRH_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH0dE+6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMD8RN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8N8sRR:#_08DHFoOC_POs0F5R4d8MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMD8RNsRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-R-RR0FsHCo#s0CRC0ERD#CCRO0#MHoNFDRVsR0HN#00NC
0H0sLCk0Rs\3NFl_VCV#0:\RRs#0H;Mo
C
Lo
HM
RRRRR--QNVR8I8sHE80RO<REOFHCH_I8R0ENH##o'MRj0'RFMRkk8#CR0LH#R
RRjRzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj"jjRN&R8C_so25j;C
SMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjjjjjjjjj"RR&Ns8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjjjjj&"RR_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjjj&"RR_N8s5CodFR8IFM0R;j2
MSC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0=ERRR62oCCMsCN0
RSRRFRDI8_N8<sR=jR"jjjjjjjj"RR&Ns8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"jjjjjjRj"&8RN_osC586RF0IMF2Rj;C
SMo8RCsMCNR0Cz
6;RRRRzRnR:VRHR85N8HsI8R0E=2R(RMoCC0sNCR
SRDRRFNI_8R8s<"=Rjjjjj"jjRN&R8C_soR5n8MFI0jFR2S;
CRM8oCCMsCN0R;zn
RRRRRz(RH:RVNR58I8sHE80RU=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjj"jjRN&R8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FINs88RR<="jjjjRj"&8RN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FINs88RR<="jjjj&"RR_N8s5CogFR8IFM0R;j2
MSC8CRoMNCs0zCRgR;
RzRR4RjR:VRHR85N8HsI8R0E=4R42CRoMNCs0SC
RRRRD_FINs88RR<="jjj"RR&Ns8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8N8s=R<Rj"j"RR&Ns8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8N8s=R<R''jRN&R8C_so.54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz.R;
RzRR4RdR:VRHR85N8HsI8R0E>dR42CRoMNCs0SC
RRRRD_FINs88RR<=Ns8_C4o5dFR8IFM0R;j2
MSC8CRoMNCs0zCR4
d;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzR4cRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rcz4;R
RR4Rz6:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
MSC8CRoMNCs0zCR4
6;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRR4RnR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s2CoRoLCHRM
RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0CRM
RRRRRRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRR(z4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_CIo5HE80-84RF0IMF2Rj;C
SMo8RCsMCNR0Cz;4(
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRp-i
-RRRRnz4RRR:H5VRNs88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCH-M
-RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Cz;4n
R--RzRR4:(RRRHV50MFR8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRNs8_C<oR=7Rq7
);-C-SMo8RCsMCNR0Cz;4(
RSRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>cR4Ro2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FRc<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;c2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.j:VRHR85N8HsI8R0E>cR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FRc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMFcR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
j;SR--Q5VRNs88I0H8E=R<R24cRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4z.RH:RVNR58I8sHE80RR<=4Rc2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vn_4dXUc4RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vn_4dXUc4RR:)Aqv41n_4R
SRRRRRRRRRbRRFRs0lRNb557Qj=2R>MRH_osC5,[2R7q7)>R=RIDF_8N8sd54RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57mj=2R>kRF0k_L#H45,2[2;R
RRRRRRRRRRRRRRkRF0C_so25[RR<=F_k0L4k#5[H,2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R.z.;R
RRSRRCRM8oCCMsCN0Rgz4;R
RRMRC8CRoMNCs0zCR4RU;R
RRRRRRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNCS
S-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzE:	RRRHV58RN8HsI8R0E>dR42CRoMNCs0RC
RRRRRzRRO:D	RFbsO#C#Rp5BiS2
RRRRRCRLo
HMSRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
SRRRRRRRRRsN8CNo58I8sHE80-84RF0IMFdR42=R<R_N8s5CoNs88I0H8ER-48MFI04FRd
2;SRSRR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5sN8CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.RX.:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qvU.4gX:.RRv)qA_4n1S.
RRRRRRRRRRRRb0FsRblNRQ57RR=>HsM_C.o5*4[+RI8FMR0F.2*[,7Rq7=)R>FRDI8_N84s5.FR8IFM0R,j2RR h='>R4R',1R1)='>RjR',
SSSSRW =I>RsC0_M25H,pRBi>R=RiBp,mR75R42=F>RkL0_k5#.H*,.[2+4,mR75Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CS-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRz	OERH:RVNR58I8sHE80R4>R.o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR.<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;.2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnXRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gcjnRXc:qR)vnA4_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Coc+*[dFR8IFM0R[c*2q,R7R7)=D>RFNI_858s484RF0IMF2Rj,hR RR=>',4'R)11RR=>',j'RS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25dRR=>F_k0Lck#5RH,c+*[dR2,7.m52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSS57m4=2R>kRF0k_L#Hc5,[c*+,42R57mj=2R>kRF0k_L#Hc5,*Rc[;22
RRRRRRRRRRRRRRRR0Fk_osC5[c*2=R<R0Fk_#Lkc,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+4RR<=F_k0Lck#5cH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*.[+2=R<R0Fk_#Lkc,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[d<2R=kRF0k_L#Hc5,[c*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
.;RRRRRMSC8CRoMNCs0zCR.
g;RRRRCRM8oCCMsCN0RUz.;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAng_1
dSzdRR:H5VROHEFOIC_HE80Rg=R2CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>R4o2RCsMCN
0CRRRRRRRRz	OD:sRbF#OC#BR5p
i2SRRRRLRRCMoH
RSRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CSM
RRRRRRRRR8RNs5CoNs88I0H8ER-48MFI04FR4<2R=8RN_osC58N8s8IH04E-RI8FMR0F4;42
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSczdRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R42M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRd6:VRHR85N8HsI8R0E>4R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF4R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
6;SR--Q5VRNs88I0H8E=R<R244RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnzdRH:RVNR58I8sHE80RR<=4R42oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_.cUUXRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_c.jURXU:qR)vnA4_
1gSRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7R7)=D>RFNI_858s48jRF0IMF2Rj,hR RR=>',4'R)11RR=>',j'RS
SS SWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm25(RR=>F_k0LUk#5UH,*([+27,Rm25nRR=>F_k0LUk#5UH,*n[+2
,RSSSS76m52>R=R0Fk_#LkU,5HU+*[6R2,7cm52>R=R0Fk_#LkU,5HU+*[cR2,7dm52>R=R0Fk_#LkU,5HU+*[dR2,
SSSS57m.=2R>kRF0k_L#HU5,[U*+,.2R57m4=2R>kRF0k_L#HU5,[U*+,42R57mj=2R>kRF0k_L#HU5,[U*2
,RSSSS75Quj=2R>MRH_osC5[g*+,U2Ru7m5Rj2=b>RN0sH$k_L#HU5,2[2;R
RRRRRRRRRRRRRRkRF0C_so*5g[<2R=kRF0k_L#HU5,[U*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*4[+2=R<R0Fk_#LkU,5HU+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[.<2R=kRF0k_L#HU5,[U*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rd2<F=RkL0_k5#UH*,U[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+cRR<=F_k0LUk#5UH,*c[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*6[+2=R<R0Fk_#LkU,5HU+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[n<2R=kRF0k_L#HU5,[U*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R(2<F=RkL0_k5#UH*,U[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+URR<=bHNs0L$_k5#UH[,R2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRSRRCRM8oCCMsCN0R(zd;R
RRSRRCRM8oCCMsCN0Rczd;R
RRMRC8CRoMNCs0zCRd
d;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n1
4USUzdRH:RVOR5EOFHCH_I8R0E=UR42CRoMNCs0SC
SR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHRN5R8I8sHE80R4>RjRR2oCCMsCN0
RRRRRRRRDzO	b:RsCFO#5#RB2pi
RSRRRRRLHCoMR
SRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRRRRRRRRNRR8osC58N8s8IH04E-RI8FMR0F4Rj2<N=R8C_so85N8HsI8-0E4FR8IFM0R24j;S
SRCRRMH8RVS;
S8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMNR58osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM5_N8s5CoNs88I0H8ER-48MFI04FRj=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;cj
-S-RRQV58N8s8IH0<ER=jR42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRcSz4RR:H5VRNs88I0H8E=R<R24jRMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;c4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRc.:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_jX.c4:nRRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq4v_jX.c4:nRRv)qA_4n1
4USRRRRRRRRRRRRsbF0NRlb7R5Q>R=R_HMs5Co4[U*+R468MFI04FRU2*[,7Rq7=)R>FRDI8_N8gs5RI8FMR0FjR2, =hR>4R''1,R1=)R>jR''
,RSSSSW= R>sRI0M_C5,H2RiBpRR=>B,piR57m4R62=F>RkL0_kn#454H,n+*[4,62R57m4Rc2=F>RkL0_kn#454H,n+*[4,c2RS
SSmS7524dRR=>F_k0L4k#n,5H4[n*+24d,mR7524.RR=>F_k0L4k#n,5H4[n*+24.,mR75244RR=>F_k0L4k#n,5H4[n*+244,SR
S7SSmj542>R=R0Fk_#Lk4Hn5,*4n[j+427,Rm25gRR=>F_k0L4k#n,5H4[n*+,g2R57mU=2R>kRF0k_L#54nHn,4*U[+2S,
S7SSm25(RR=>F_k0L4k#n,5H4[n*+,(2R57mn=2R>kRF0k_L#54nHn,4*n[+27,Rm256RR=>F_k0L4k#n,5H4[n*+,62
SSSRRRR7cm52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR75Rd2=F>RkL0_kn#454H,n+*[dR2,7.m52>R=R0Fk_#Lk4Hn5,*4n[2+.,S
SRRRRRRRR74m52>R=R0Fk_#Lk4Hn5,*4n[2+4,mR75Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7QRR=>HsM_C4o5U+*[48(RF0IMFUR4*4[+n
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u254RR=>bHNs0L$_kn#45RH,.+*[4R2,75muj=2R>NRbs$H0_#Lk4Hn5,*R.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRc
.;RRRRRMSC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nz
Sc:dRRRHV5FOEH_OCI0H8ERR=dRn2oCCMsCN0
-SS-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRR8N8s8IH0>ERR2gRRMoCC0sNCR
SRzRRO:D	RFbsO#C#Rp5BiS2
SLRRCMoH
RSSRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMSRSRRRRRNC8so85N8HsI8-0E4FR8IFM0RRg2<N=R8C_so85N8HsI8-0E4FR8IFM0R;g2
RSSRMRC8VRH;S
SCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;SRRRRczcRV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>gM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOS
SS6zcRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SFSSkC0_M25HRR<='R4'IMECR85Ns5CoNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMNR58C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc
6;SR--Q5VRNs88I0H8E=R<RRg2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
SSSzRcn:VRHR85N8HsI8R0E<g=R2CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
SSSS0Is_5CMH<2R= RW;S
SS8CMRMoCC0sNCcRznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzRc(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRRRRRR)RAq6v_4d.X.RR:)Aqv41n_dRn
RRRRRRRRRRRRRRRRRbRRFRs0lRNb5R7Q=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77RD=>FNI_858sUFR8IFM0R,j2RR h='>R4R',1R1)='>Rj
',RRRRRRRRRRRRRRRRRRRRRRRRRRRRR RWRR=>I_s0CHM52B,Rp=iR>pRBi7,Rm45d2>R=R0Fk_#LkdH.5,*d.[4+d27,Rmj5d2>R=R0Fk_#LkdH.5,*d.[j+d2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rg2=F>RkL0_k.#d5dH,.+*[.,g2R57m.RU2=F>RkL0_k.#d5dH,.+*[.,U2R57m.R(2=F>RkL0_k.#d5dH,.+*[.,(2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmn5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm65.2>R=R0Fk_#LkdH.5,*d.[6+.27,Rmc5.2>R=R0Fk_#LkdH.5,*d.[c+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.Rd2=F>RkL0_k.#d5dH,.+*[.,d2R57m.R.2=F>RkL0_k.#d5dH,.+*[.,.2R57m.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmj5.2>R=R0Fk_#LkdH.5,*d.[j+.27,Rmg542>R=R0Fk_#LkdH.5,*d.[g+427,RmU542>R=R0Fk_#LkdH.5,*d.[U+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m4R(2=F>RkL0_k.#d5dH,.+*[4,(2R57m4Rn2=F>RkL0_k.#d5dH,.+*[4,n2R57m4R62=F>RkL0_k.#d5dH,.+*[4,62
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmc542>R=R0Fk_#LkdH.5,*d.[c+427,Rmd542>R=R0Fk_#LkdH.5,*d.[d+427,Rm.542>R=R0Fk_#LkdH.5,*d.[.+42
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR75244RR=>F_k0Ldk#.,5Hd[.*+244,mR7524jRR=>F_k0Ldk#.,5Hd[.*+24j,mR75Rg2=F>RkL0_k.#d5dH,.+*[gR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm25URR=>F_k0Ldk#.,5Hd[.*+,U2R57m(=2R>kRF0k_L#5d.H.,d*([+27,Rm25nRR=>F_k0Ldk#.,5Hd[.*+,n2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR76m52>R=R0Fk_#LkdH.5,*d.[2+6,mR75Rc2=F>RkL0_k.#d5dH,.+*[cR2,7dm52>R=R0Fk_#LkdH.5,*d.[2+d,RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR57m.=2R>kRF0k_L#5d.H.,d*.[+27,Rm254RR=>F_k0Ldk#.,5Hd[.*+,42R57mj=2R>kRF0k_L#5d.H.,d*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RQu=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,Rmdu52>R=RsbNH_0$Ldk#.,5HR[c*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.u52>R=RsbNH_0$Ldk#.,5HR[c*+,.2Ru7m5R42=b>RN0sH$k_L#5d.Hc,R*4[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7m5Rj2=b>RN0sH$k_L#5d.Hc,R*2[2;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*4[+2=R<R0Fk_#LkdH.5,*d.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*d[+2=R<R0Fk_#LkdH.5,*d.[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*6[+2=R<R0Fk_#LkdH.5,*d.[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*([+2=R<R0Fk_#LkdH.5,*d.[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRRkRF0C_son5d*g[+2=R<R0Fk_#LkdH.5,*d.[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+244RR<=F_k0Ldk#.,5Hd[.*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24dRR<=F_k0Ldk#.,5Hd[.*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+246RR<=F_k0Ldk#.,5Hd[.*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24(RR<=F_k0Ldk#.,5Hd[.*+24(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+24gRR<=F_k0Ldk#.,5Hd[.*+24gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.4RR<=F_k0Ldk#.,5Hd[.*+2.4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.dRR<=F_k0Ldk#.,5Hd[.*+2.dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.6RR<=F_k0Ldk#.,5Hd[.*+2.6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.(RR<=F_k0Ldk#.,5Hd[.*+2.(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2.gRR<=F_k0Ldk#.,5Hd[.*+2.gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d4RR<=F_k0Ldk#.,5Hd[.*+2d4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRRFRRks0_Cdo5n+*[dRd2<b=RN0sH$k_L#5d.H*,c[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRRRRF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRRRRR0Fk_osC5*dn[6+d2=R<RsbNH_0$Ldk#.,5Hc+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SCSSMo8RCsMCNR0Cz;c(
CSSMo8RCsMCNR0Cz;cc
MSC8CRoMNCs0zCRc
d;CRM8NEsOHO0C0CksR_MFsOI_E	CO;-

--
-R#pN0lRHblDCCNM00MHFRRH#8NCVk
D0-N-
sHOE00COkRsC#CCDOs0_NFlRVqR)vW_)u#RH
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;O#FM00NMRlMk_DOCD:#RR0HMCsoCRR:=5C58bR0E-2R4/24n;RRRRRRRRRRRRR--yVRFRv)q44nX7CRODRD#M8CCC08
$RbCF_k0L_k#0C$bRRH#NNss$MR5kOl_C#DDRI8FMR0FjI,RHE80-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#RR:F_k0L_k#0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_RCM:0R#8F_Do_HOP0COFMs5kOl_C#DDRI8FMR0FjR2;RRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRR-R-RCk#8FR0RosCHC#0sQR7h#R
HNoMDkRF0C_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNR8N8s0_#oRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-b-RHDbCHRMCs8CNRosCHC#0s0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RRcNH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR8N8s0_#o25j;R
RRRRRRFRDIN_I8R8s<"=Rj"jjRN&R8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8N8s0_#oR548MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=""jjRN&R8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR8N8s0_#oR5.8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<='Rj'&8RN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0>ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=8RN8#s_0do5RI8FMR0Fj
2;RRRRRRRRD_FII8N8s=R<R_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR6RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=7;Qh
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRz(RH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
pi-R-RRgRzRRR:H5VRNs88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#Rp5Biq,R727)RoLCH-M
-RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR_N8sRCo<q=R757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-R-RRMRC8CRoMNCs0zCRg-;
-RRRRjz4RH:RVMR5FN0R8_8ss2CoRMoCC0sNCR
RRRRRRRRRR8RN_osCRR<=q)77;-
-RRRRCRM8oCCMsCN0Rjz4;R
RRRRRRRR
R-RR-HRbbHCDM#CR0CNo8CRso0H#CRs
RzRR4R6R:sRbF#OC#BR5pRi,Ns8_C
o2SRRRLHCoMR
RRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRNs88_o#0RR<=Ns8_CNo58I8sHE80-84RF0IMF2Rj;R
RRRRRRMRC8VRH;R
RRMRC8sRbF#OC#4Rz6R;
R
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHRO
RzRR4:4RRsVFRHHRMkRMlC_ODRD#8MFI0jFRRMoCC0sNCR
RRRRRR-R-RRQV58N8s8IH0>ERRRc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4:.RRRHV58N8s8IH0>ERRRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRNs88_o#058N8s8IH04E-RI8FMR0Fc=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRNs8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0R.z4;R
RRRRRR-R-RRQV58N8s8IH0<ER=2RcRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR4RzdRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRRRRRCRM8oCCMsCN0Rdz4;R
RR-R-RCtMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRR4RzcRR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzq:vRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo54H*n&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E5+HRR*424Rn,80CbER22&XR""RR&HCM0o'CsHolNC+5[4
2;RRRRRRRRRRRRLHCoMR
RRRRRRRRRR)RzqRv:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=R_HMs5Co[R2,q=jR>FRDIN_I858sjR2,q=4R>FRDIN_I858s4R2,q=.R>FRDIN_I858s.
2,RRRRRRRRRRRRRRRRRRRRRRRRRdRqRR=>D_FII8N8s25d,uR7)Rqj=D>RFsI_Ns885,j2R)7uq=4R>FRDIN_s858s4R2,
RRRRRRRRRRRRRRRRRRRRRRRR7RRu.)qRR=>D_FIs8N8s25.,uR7)Rqd=D>RFsI_Ns885,d2RRW =I>RsC0_M25H,RR
RRRRRRRRRRRRRRRRRRRRRRRRRpWBi>R=RiBp,uR7m>R=R0Fk_#Lk5[H,2
2;RRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRCRM8oCCMsCN0Rcz4;R
RRRRRRMRC8CRoMNCs0zCR4
4;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRM
C8sRNO0EHCkO0s#CRCODC0N_sl
;

