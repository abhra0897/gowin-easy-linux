@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ha_me_m p)wm;W"
R
R`OHMDCk8R0"#8P_FDN_0#E	3"


`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vt`

HCV8VeRmp1_q1a )_
mh
bRRsCFbsR0$q 11)ha_me_m p)wmuW_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5#0C0G_Cb=sR=NRlG|2R=5>R5#0C0G_Cb>sRRMlH2&R&RC50#C0_GRbs<l=RN2G2;R
RCbM8sCFbs
0$R
R
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
bRRsCFbsR0$q 11)ha_me_m p)wmXW_Zh_m_1a aX_ uu)_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5HM#k	IMFMC50#C0_G2bs2
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRR_Rqq 11)ha_me_m p)wmuW_:#RN#0CsRFbsb0Cs$qR51)1 am_h_ me)mwpW2_u
RRRRRRRR#CDCPRFDs_Cs_Fs0a5"CR#0CsGbCH##FOMREoNMCP8RNCDkRFVslDRNDCFI8NRlGkHllNRPDRkClRNG0NFRRDPNkHCRMER0CNRsMRoCl+NG4FR0RMlH"
2;
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRqRR_1q1 _)ahmm_ew )p_mWXmZ_h _a1 a_X_u)uR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)ha_me_m p)wmXW_Zh_m_1a aX_ uu)_2R
RRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2RRR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w

RRRRCRRMR8
RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRR_Rvq 11)ha_me_m p)wmuW_:#RN#CklRFbsb0Cs$qR51)1 am_h_ me)mwpW2_u;`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )__hmm)e wWpm__XZmah_ _1a )Xu_
u:RRRRRRRRNk##lbCRsCFbsR0$51q1 _)ahmm_ew )p_mWXmZ_h _a1 a_X_u)uR2;
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR7R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
R
RRVRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRRRH5VRm_epB me)q_A1_QBmRh2LHCoMRR:F_PDOCFPsN_L#
HORRRRRR
RRRRROCFPsC_0#C0_G_bsNl0_N
G:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRf#sFCC50#C0_GRbs=l=RNRG22R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbNs_0N_lGFROPCCs8;"2
RRRRMRC8/R/LHN#OFROPNCso
C
RRRRRRHV5pme_eBm B)_m )h)h_m2CRLoRHM:PRFDF_OP_CsOMFsC
s
RRRRRFROP_Cs00C#_bCGs0_N_MlH:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRsRfF5#C00C#_bCGs=R=RMlH22R2
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb__N0lRHMOCFPs"C82R;
RRRRCRM8/F/OssMCRPOFCosNCR
RRMRC8C

MC8oMNCs0
C
`8CMH/VR/eRmpm_Be_ )m
h

