-- --------------------------------------------------------------------
@E
---B-RFsb$H0oER.�RjRjULQ$R 3  RDqDRosHER0#sCC#s8PC3-
-
R--a#EHRk#FsROCVCHDRRH#NCMR#M#C0DHNRsbN0VRFR Q  0R18jR4(.n-j,jU
R--Q   RN10Ms8N8]Re7ppRNkMoNRoC)CCVsOCMCNRvMDkN3ERaH##RFOksCHRVDlCRNM$RFL0RC-
-RbOFH,C8RD#F8F,RsMRHO8DkCI8RHR0E#0FVICNsRN0E0#RHRD#F8HRI0kEF0sRIHC00M-R
-CRbs#lH#MHFRFVslER0C RQ 1 R08NMN#s8Rb7CNls0C3M0RHaE#FR#kCsORDVHCNRl$CRLR-
-RbOFHRC8VRFsHHM8PkH8NkDR#LCRCC0ICDMRHMOC#RC8ks#C#a3RERH##sFkOVCRHRDCH-#
-sRbF8PHCF8RMMRNRRq1QL1RN##H3ERaC RQ 8 RHD#ON#HlRYqhR)Wq)aqhYXR u1) 1)Rm
R--QpvuQR 7QphBzh7QthRqYqRW)h)qamYRw Rv)qB]hAaqQapQYhRq7QRwa1h 1mRw)1Rz -
-R)wmRuqRqQ)aBqzp)zRu)1um a3REkCR#RCsF0VRE#CRFOksCHRVD#CREDNDR8HMCHlMV-$
-MRN8FREDQ8R R  ElNsD#C#RFVslMRN$NR8lCNo#sRFRNDHLHHD0N$RsHH#MFoRkF0RVER0C-
-RCk#RC0EsVCF3-
-
R--RHRa0RDCRRRR:wRRD0FNH-MobMFH0NRbOo	NCQR5MN#0MN0H0RC8b	NONRoC8DCON0sNH2FM
R--RRRRRRRRRRRR:-
-RpRRHNLssR$RRR:Ra#EHRObN	CNoRN#EDLDRCFROlDbHCH8RMR0FNHRDLssN$-
-RRRRRRRRRRRRRR:R#L$lFODHN$DDRlMNCQ8R 3  
R--RRRRRRRRRRRR:-
-R7RRCDPCFsbC#R:RqCOODsDCN]Re7ap-BMRN8 RQ u R4nj(RsWF	oHMRFtsk-b
-RRRRRRRRRRRR
R:-R-RRsukbCF#R:RRRERaHb#RNNO	oRC#8HCVMRC#LHN#OHRLM$NsRFVDNM0HoFRbH
M0-R-RRRRRRRRRR:RRRsRNHl0ECO0HRMVkOF0HM-#
-RRRRRRRRRRRR
R:-R-RR0hFCRRRR:RRRERaHb#RNNO	olCRNL$RCFRl8HHVC08RFMRHO8DkC8RN8HH0FDMNR08NN-
-RRRRRRRRRRRRRR:RskCJH8sCRRL$0DFF#L,RkH0R0kRl#H0RMFRMR$INRNOEMRoC0
EC-R-RRRRRRRRRR:RRRGRC0MCsNHDRMs0CVCNO#sRFRl#Hk0DNHRFMLNCEPsHFRRFV0
EC-R-RRRRRRRRRR:RRRCR8#HOsbF0HMQ3R0#RHRsbCl#H#HCLDRR0FNR88OlFlC#M0R8NM/
Fs-R-RRRRRRRRRR:RRR0RN0LsHk#0CRR0F0RECb	NONRoC8DCON0sNH#FM,kRL0FRM0FR0RNOEM
oC-R-RRRRRRRRRR:RRRsRFRD8CCR0CNRM$FosHHDMNRMDHCF#RVER0CNRbOo	NCCR8OsDNNF0HM-3
-RRRRRRRRRRRRRR:RCaERObN	CNoR8LF$NRl$CRLRNOEM8oCRDFM$MRHRONOFNs8MROCIEH0
R--RRRRRRRRRRRR:0RRE0CRC#slRRFVBkDN#4CRnVRFRH0E#0R#NNM8s
83-R-RRRRRRRRRR:RR
R----------------------------------------------------------------------
R--fP)CHF#HM4:R.R.jf-
-RNf70RC:.Ujj--jc44jR(n:4:Rjg+djgjaR5ERk,4qjRb.sRj2jUR-f
--R------------------------------------------------------------------
-
DsHLNRs$HCCC;b

NNO	oVCRD0FN_ob	RRH#MRCIQ   3FVDNo0_CsMCHbO_	Ro
RMoCCOsHRblNRR5
RVRRD0FN_ksFM#8_0C$DRRRR=Q>R 3  VCHG8D_VF_N00C$b#F3sk_M8MsCNC,#0R-R-RksFMM8RCCNs#N0RDsoFHl0E
RRRRFVDNC0_GMbFC_M0I0H8E>R=RRU,R-RR-DRVFdN0.H'EoRE
RVRRD0FN_NVsOF0HMH_I8R0E=.>RdR,RRR---FVDN.0d'IDF
RRRRFVDN80_CsMFlHNDxRCRR>R=Rk0sCR,R-z-R#QCR R  CCG0M88CRFVDNM0HoR
RRDRVF_N0OOEC	s_CsRFsR=RR>sR0kRC,RR--aMksRRFMhRqhNRM8FsPCVIDFRFbsO#C#H
MoRRRRVNDF0k_oN_s8L#H0RRRRRR=>dR,RR-RR-kRMlsLCRRFVoskN8HRL0R#
RMRRFN_IsMMHoRRRRRRRRRRR=V>RNCD#RR--#IEFRsINMoHM#R
RR;R2
