@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)a7) B hv a
";
V`H8RCVm_epQahQ_tv1
HRRMHH0NRD
RFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8
HV
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_B7 )  vhua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5#L0ND0C5C_#0CsGb2&2R&bRfN5#0`pme_1)  1a_Qqthp22RR>|-R55R00C#_bCGsRR<f#bN0C50#C0_G2bs2
R?RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RRf#bN0C50#C0_G2bsR0-RC_#0CsGbRR==PkNDC:2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5Nfb#005C_#0CsGb2RR+5H{I8{0E44'L}-}RR#0C0G_CbRs2+'R4L=4R=NRPD2kC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2R;
R8CMbbsFC$s0
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRsRbFsbC0q$R1)1 a _7Bv)  _haXmZ_h _a1 a_X_u)uR;
RR@@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )_B7 )  vhua_:R
RRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _7Bv)  _hauC2RDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRRH#8sCOCCN#8$RLRPNRNCDkREF0C0sRERNM#ObCHCVH8;"2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRqRR_1q1 _)a7) B hv aZ_X__mhaa 1_u X):_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_B7 )  vhXa_Zh_m_1a aX_ uu)_2R
RRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRM
8
RRRRRmR`eqp_1v1z RR:LHCoMRR:F_PDNk##lRC
RRRRRvRR_1q1 _)a7) B hv a:_uR#N#kRlCbbsFC$s0R15q1a )_B7 )  vhua_2
;R
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rvq 11)7a_  B)va h__XZmah_ _1a )Xu_
u:RRRRRRRRNk##lbCRsCFbsR0$51q1 _)a7) B hv aZ_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
RCRoMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RRRRRPOFC0s_C_#0CsGb_NOEM:oC
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR!RRfN#0L5DC00C#_bCGs22R2R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsE_ONCMoRPOFC8sC"
2;RRRRR8CM
RRRR8CM
R
RCoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
