@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)za_hqB]h"t ;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"
`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vtR

RHHM0DHNRoLCHRM
RHRRV5R5M_klOR	#<2=jR
||RRRRRRRR~N55OF0HMM_F_IMC_N#0s=0R=mR`eQp_t)hm  _hWa_1q2)aR
||RRRRRRRRRNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqa|2R|R
RRRRRRRRR50NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)a2L2RCMoH
RRRRFRRPCD_sssF_"05QCDDoRNDPkNDCCR#0FRVsNRbsCNl0RCsNHO0FFM_MC_MI0_#NRs0FbsRNlsNCs0CRlMk_#O	"
2;RRRRC
M8RMRC8
RR
V`H8RCVm_ep1)]q B7_m
7 
sRRCIoRHFM8IRR=jR;
R0HMCsoCR=HRR
j;
NRRD$IN#@R@RF5b#oC8CDRO	L2RCMoH
RRRRRHV5e`mp _)1_ a1hQtq!pR='R4LRj2LHCoMR
RRRRRH5VR!MIH8RFI&#&R00Ns_CCPM=0R='R4LR42LHCoMR
RRRRRRHRIMI8FRR<=44'L;R
RRRRRRRRH<M=RkOl_	
#;RRRRRMRC8R
RRRRRCCD#RRHV5MIH82FIRoLCHRM
RRRRRHRRVHR5RR==4&R&RO5N0MHF__FMM_CI#s0N0=R!Re`mp _)1_ amhh_ 1W_aaq)RR||#s0N0P_CCRM0!4=R'2L42R
RRRRRRRRRI8HMF<IR='R4L
j;
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_1)  ma_h _hWa_1qR)a&#&R00Ns_CCPM=0R='R4L
42RRRRRRRRRRRH<M=RkOl_	
#;RRRRRRRRCCD#RRHV5!HR=2R4
RRRRRRRRHRRRR<=HRR-4R;
RRRRR8CMRR//H5VRI8HMF
I2RRRRC
M8RRRRCCD#RoLCHRM
RRRRRMIH8RFI<4=R';Lj
RRRRHRRRR<=jR;
RCRRMR8
R8CM
C
`MV8HRR//m_ep1)]q B7_m
7 
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_Bzh]tqh ;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RR#s0N0P_CCRM0&!&RI8HMFRI2|R=>50f#NCLD5#0C0G_Cbrs2*lMk_#O	9
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_Bzh]tqh  _)1_ am1h_aaq)_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R#R500Ns_CCPMR02|R=>5RR
RRRRRRRRRRRRRRRRRRRRR#5f0DNLCC50#C0_G2bsrk*Ml	_O#
92SRRRRRRRRRRRRFRRsRR
RRRRRRRRRRRRRRRRRRRRR#5f0DNLCC50#C0_G2bsr:*jM_klO-	#4y9Ry#4R00Ns_CCPMR02
RSRRRRRRRRRR;R2
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 ah_zBh]qt  _)m)_ha_1q_)auR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RMIH8RFI|R->!N#0sC0_P0CM;R
RCbM8sCFbs
0$
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RbbsFC$s0R1q1 _)az]hBq ht__XZm1h_aaq)_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R!I8HMFRI2|R->5f!5HM#k	IMFM05#N_s0CMPC0222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)za_hqB]h_t XmZ_h _hWa_1q_)auR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RH5IMI8F2-R|>!R55#fHkMM	F5IM#s0N0P_CC2M02
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_Bzh]tqh Z_X__mhaa 1_u X);_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRI8HMF|IR|0R#N_s0CMPC0|2R-5>R!H5f#	kMMMFI5#0C0G_Cb2s22R;
R8CMbbsFC$s0
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
oRRCsMCN
0CRRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_ep)  1ah_m_Wh _q1a)
a2RRRRRRRRR_Rqq 11)za_hqB]h_t uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Bzh]tqh 2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRNOEM8oCRDPNkICRHH0EMkRMl	_O#sRVF0lRE#CR00NsRCCPMN0R#s#C0"C82R;
RRRRRHRRVNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqaR2
RRRRRRRRRqq_1)1 ah_zBh]qt) _ a1 __mh1)aqa:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)za_hqB]h_t )  1ah_m_q1a)ua_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HMERONCMo8NRPDRkCIEH0HMMRkOl_	V#RsRFl0REC#s0N0PRCCRM0NC##s80C"
2;RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0=`=Rm_ep m)))h_m_Wh _q1a)
a2RRRRRRRRR_Rqq 11)za_hqB]h_t  _))m1h_aaq)_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ah_zBh]qt  _)m)_ha_1q_)auR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0Q5"DoDCN#DR00NsRCCPMI0REEHOR#ENRFsCOsOkCL8RCsVFCFROlCbD0MHFRRFVOsksCRM0I8HMF2I";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRRRRq1_q1a )_Bzh]tqh Z_X__mh1)aqa:_u
RRRRRRRRRRRNC##sb0RsCFbsR0$51q1 _)az]hBq ht__XZm1h_aaq)_
u2RRRRRRRRRCRRDR#CF_PDCFsss5_0"N#0sC0_P0CMRMOF0MNH#RRXFZsR"
2;RRRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR!=`pme_hQtm_) h_ W1)aqaR2
RRRRRRRRR_Rqq 11)za_hqB]h_t XmZ_h _hWa_1q_)auR:
RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ah_zBh]qtX _Zh_m_Wh _q1a)ua_2R
RRRRRRRRRR#CDCPRFDs_Cs_Fs0#5"00Ns_CCPMO0RFNM0HRM#XsRFR2Z";R
RRRRRRqRR_1q1 _)az]hBq ht__XZmah_ _1a )Xu_
u:RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Bzh]tqh Z_X__mhaa 1_u X)2_u
RRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R!Re`mp _)1_ amhh_ 1W_aaq)2R
RRRRRRRRRv1_q1a )_Bzh]tqh :_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)za_hqB]h_t u
2;RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0=`=Rm_ep)  1ah_m_Wh _q1a)
a2RRRRRRRRR_Rvq 11)za_hqB]h_t )  1ah_m_q1a)ua_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)az]hBq ht_1)  ma_ha_1q_)au
2;RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0=`=Rm_ep m)))h_m_Wh _q1a)
a2RRRRRRRRR_Rvq 11)za_hqB]h_t  _))m1h_aaq)_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 ah_zBh]qt  _)m)_ha_1q_)au
2;
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRRRRR_Rvq 11)za_hqB]h_t XmZ_ha_1q_)auR:
RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 ah_zBh]qtX _Zh_m_q1a)ua_2R;
RRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_epQmth)h _ 1W_aaq)2R
RRRRRRRRRRqv_1)1 ah_zBh]qtX _Zh_m_Wh _q1a)ua_:R
RRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Bzh]tqh Z_X__mhh_ W1)aqa2_u;R
RRRRRRvRR_1q1 _)az]hBq ht__XZmah_ _1a )Xu_
u:RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Bzh]tqh Z_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_ho

CsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_CsI8HMFFI_b:CM
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRRRRRN#0sC0_P0CMRR&&!MIH82FIRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8_FIFMbCRPOFC8sC"
2;
RRRRORRFsPC_MIH8_FIO#DFCR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRRRRRRRRRRRRRRIRRHFM8I&R&RR5H=4=RRR&&50NOH_FMFMM_C#I_00NsRR!=`pme_1)  ma_h _hWa_1qR)a|#|R00Ns_CCPM!0R='R4L2422
R2RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5H"IMI8F_FOD#OCRFsPCC28";R
RRCRRM/8R/#LNHOORFsPCN
oC
RRRRVRHRe5mpm_Be_ )Bhm) m)_hL2RCMoHRF:RPOD_FsPC_sOFM
CsRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2CRLoRHM:PRFDF_OP_CsI8HMFsI_C0#C#R
RRRR
RRRRRFROP_CsI8HMFsI_C0#C#R:
RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRR#s0N0P_CCRM0&I&RHFM8I22R
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs0I5"HFM8IC_s##C0RPOFC8sC"
2;RRRRRMRC8R
RRCRRM/8R/sOFMRCsOCFPsCNo
RRRR8CM
M
C8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



