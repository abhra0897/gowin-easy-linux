@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)qa_pYWq1h_m_t 7 
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E

RR`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vt`

HCV8VeRmp1_q1a )_
mh
bRRsCFbsR0$q 11)qa_pYWq1h_m_t 7 m_h  7t_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RCR0#C0_G;bs
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_1um  7t_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RyR5yf4RsCF#5l#NbMDHoP_CC2M02-R|>CR0#C0_G;bs
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_th   7t_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RyR5yf4RVDCD5l#NbMDHoP_CC2M02-R|>CR0#C0_G;bs
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_Yqh  7t_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RyR5y!4R50f#NCLD5l#NbMDHoP_CC2M02|2R-0>RC_#0CsGb;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RbRRsCFbsR0$q 11)qa_pYWq1h_m_t 7 m_h  7t_1a aX_ uX)_Z;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRRf5!HM#k	IMFMC50#C0_G2bs2R;
RCRRMs8bFsbC0
$
RRRRbbsFC$s0R1q1 _)aqqpWYm1_h7_ tu _m71 t1 _q_vu he a__jXuZ_;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RR5R5yRy45!R5f#bN0N5#lHbDMCo_P0CM2222R>|-Rf5!HM#k	IMFMN5#lHbDMCo_P0CM2;22
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_1um  7t_v1que_  _haX4Z__
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5y5y45R5fkH#MF	MIfM5b0N#5l#NbMDHoP_CC2M02&2R&!R5fkH#MF	MI#M5NDlbH_MoCMPC02222R
RRRRR|R->5N!#lHbDMCo_P0CM2
2;RRRRCbM8sCFbs
0$
RRRRFbsb0Cs$1Rq1a )_Wqpq_Y1m h_7_t 1uqv_  ehXa_ZZ_X_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5yR5yR4R5#fHkMM	F5IM#bNlDoHM_CCPM2022RR
RRRRR>|-Rf5!HM#k	IMFMb5fN5#0#bNlDoHM_CCPM2022;R2
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_1um  7t_1a aX_ uX)_Z;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRRy55yf4RsCF#5l#NbMDHoP_CC2M02-R|>!R5fkH#MF	MI0M5C_#0CsGb2;22
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_th   7t_v1que_  _ha4Z_X_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5yR5y54Rf#bN0N5#lHbDMCo_P0CM2R22|R->5H!f#	kMMMFI5l#NbMDHoP_CC2M02;R2
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_th   7t_v1que_  _haXjZ__
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5yR5y54R5#fHkMM	F5IMf#bN0N5#lHbDMCo_P0CM2222R5&&!#fHkMM	F5IM#bNlDoHM_CCPM2022R
RR|RR-5>R#bNlDoHM_CCPMR022R;
RCRRMs8bFsbC0
$
RRRRbbsFC$s0R1q1 _)aqqpWYm1_h7_ th _ 7t ta _ _1a )Xu__XZuR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R5RR54yyRCfVD#D5NDlbH_MoCMPC0R22|R->5H!f#	kMMMFI5#0C0G_Cb2s22R;
RCRRMs8bFsbC0
$
RRRRbbsFC$s0R1q1 _)aqqpWYm1_h7_ tq _h7Y t1 _q_vu he aZ_X_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5f!5HM#k	IMFMN5#lHbDMCo_P0CM2;22
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_Yqh  7t_ u)eq_1v u_ea h__XZuR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R5RRRy5y4H5f#	kMMMFI5Nfb##05NDlbH_MoCMPC02222-R|>fR5HM#k	IMFMN5#lHbDMCo_P0CM2;22
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 ap_qW1qY__mh  7t_Yqh  7t_1a aX_ uX)_Z;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRRy55y!4R50f#NCLD5l#NbMDHoP_CC2M02|2R-5>R!#fHkMM	F5IM00C#_bCGs222;R
RRMRC8Fbsb0Cs$R

RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRCC8o_b0$C=R=Re`mpm_h  7t2CRLoRHM:_RNNC##sN0_D$IN#M_F_oC8CF_MCC8o
RRRRRRRRqRR_1q1 _)aqqpWYm1_h7_ th _mt 7 :_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)qa_pYWq1h_m_t 7 m_h  7t_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHw#Rq p1RsHsCC#bOP0HCVRFRl#NbMDHoPRCC"M02
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRRRRRq1_q1a )_Wqpq_Y1m h_7_t h7m ta _ _1a )Xu__XZuR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Wqpq_Y1m h_7_t h7m ta _ _1a )Xu__XZuR2
RRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w

RRRRRRRR8CM
R
RRRRRRVRHR85Co0C_$RbC=`=Rm_epu m172t RoLCH:MRRNN_#s#C0D_NI#N$__FMCC8o_#bFCC8o
RRRRRRRRqRR_1q1 _)aqqpWYm1_h7_ tu _m71 tu _:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aqqpWYm1_h7_ tu _m71 tu _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHRpwq1F RMFRb#oC8CVRFRl#NbMDHoPRCC"M02
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRRRRRq1_q1a )_Wqpq_Y1m h_7_t u m17_t aa 1_u X)Z_X_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_1um  7t_1a aX_ uX)_Z2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"#0C0G_CbOsRFNM0HRM#XsRFR2Z";R

RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_1um  7t_v1que_  _hajZ_X_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_1um  7t_v1que_  _hajZ_X_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#bNlDoHM_CCPMO0RFNM0HRM#XsRFR2Z";R

RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_1um  7t_v1que_  _haX4Z__
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_1um  7t_v1que_  _haX4Z__
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#bNlDoHM_CCPMO0RFNM0HRM#XsRFR2Z";R

RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_v1que_  _haXXZ_Z:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)qa_pYWq1h_m_t 7 q_1v u_ea h__XZXuZ_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5N"#lHbDMCo_P0CMRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w

RRRRRRRR8CM
R
RRRRRRVRHR85Co0C_$RbC=`=Rm_eph  t72t RoLCH:MRRNN_#s#C0D_NI#N$__FMCC8o_oMCCC8o
RRRRRRRRqRR_1q1 _)aqqpWYm1_h7_ th _ 7t tu _:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aqqpWYm1_h7_ th _ 7t tu _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHRpwq1F RMCRMooC8CVRFRl#NbMDHoPRCC"M02
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRRRRRq1_q1a )_Wqpq_Y1m h_7_t h  t7_t aa 1_u X)Z_X_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_th   7t_1a aX_ uX)_Z2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"#0C0G_CbOsRFNM0HRM#XsRFR2Z";R

RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_th   7t_v1que_  _ha4Z_X_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_th   7t_v1que_  _ha4Z_X_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#bNlDoHM_CCPMO0RFNM0HRM#XsRFR2Z";R

RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_th   7t_v1que_  _haXjZ__
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_th   7t_v1que_  _haXjZ__
u2RRRRRRRRRDRC#FCRPCD_sssF_"05Rl#NbMDHoP_CCRM0O0FMN#HMRFXRsRRZ"
2;
RRRRRRRRqRR_1q1 _)aqqpWYm1_h7_ t1 _q_vu he aZ_X__XZuR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Wqpq_Y1m h_7_t 1uqv_  ehXa_ZZ_X_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05#bNlDoHM_CCPMO0RFNM0HRM#XsRFR2Z";R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R

RRRRRCRRM
8
RRRRRRRRH5VRCC8o_b0$C=R=Re`mph_qYt 7 L2RCMoHRN:R_#N#C_s0NNDI$F#_M8_CoNC_M8$CoRC
RRRRRRRRRqq_1)1 ap_qW1qY__mh  7t_Yqh  7t_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_Yqh  7t_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHw#Rq p1RRFMNRM$CC8oRRFV#bNlDoHMRCCPM20";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqRR_1q1 _)aqqpWYm1_h7_ tq _h7Y ta _ _1a )Xu__XZuR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Wqpq_Y1m h_7_t q hY7_t aa 1_u X)Z_X_
u2RRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
R
RRRRRRRRRq1_q1a )_Wqpq_Y1m h_7_t q hY7_t 1uqv_  ehXa_Z:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)qa_pYWq1h_m_t 7 h_qYt 7 q_1v u_ea h__XZuR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0#5"NDlbH_MoCMPC0FROMH0NMX#RRRFsZ;"2
R
RRRRRRRRRq1_q1a )_Wqpq_Y1m h_7_t q hY7_t ue) _v1que_  _haXuZ_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aqqpWYm1_h7_ tq _h7Y tu _)_ e1uqv_  ehXa_Z2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"l#NbMDHoP_CCRM0O0FMN#HMRFXRs"RZ2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRC
M8RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRRHV5oC8C$_0b=CR=mR`ehp_mt 7 L2RCMoHRl:R_#N#C_s0NNDI$F#_M8_CoMC_FoC8CR
RRRRRRRRRv1_q1a )_Wqpq_Y1m h_7_t h7m tu _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aqqpWYm1_h7_ th _mt 7 2_u;


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRvRR_1q1 _)aqqpWYm1_h7_ th _mt 7  _a1 a_X_u)XuZ_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aqqpWYm1_h7_ th _mt 7  _a1 a_X_u)XuZ_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRC
M8
RRRRRRRRRHV5oC8C$_0b=CR=mR`eup_m71 tR 2LHCoMRR:l#_N#0Cs_INDN_$#FCM_8_oCbCF#8
oCRRRRRRRRR_Rvq 11)qa_pYWq1h_m_t 7 m_u1t 7 :_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)qa_pYWq1h_m_t 7 m_u1t 7 2_u;


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRvRR_1q1 _)aqqpWYm1_h7_ tu _m71 ta _ _1a )Xu__XZuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t u m17_t aa 1_u X)Z_X_;u2
R
RRRRRRRRRv1_q1a )_Wqpq_Y1m h_7_t u m17_t 1uqv_  ehja___XZuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t u m17_t 1uqv_  ehja___XZu
2;
RRRRRRRRvRR_1q1 _)aqqpWYm1_h7_ tu _m71 t1 _q_vu he aZ_X_u4_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aqqpWYm1_h7_ tu _m71 t1 _q_vu he aZ_X_u4_2
;
RRRRRRRRR_Rvq 11)qa_pYWq1h_m_t 7 q_1v u_ea h__XZXuZ_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aqqpWYm1_h7_ t1 _q_vu he aZ_X__XZu
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w

RRRRRRRR8CM
R
RRRRRRVRHR85Co0C_$RbC=`=Rm_eph  t72t RoLCH:MRRNl_#s#C0D_NI#N$__FMCC8o_oMCCC8o
RRRRRRRRvRR_1q1 _)aqqpWYm1_h7_ th _ 7t tu _:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aqqpWYm1_h7_ th _ 7t tu _2
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRRRRRv1_q1a )_Wqpq_Y1m h_7_t h  t7_t aa 1_u X)Z_X_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_th   7t_1a aX_ uX)_Z2_u;R

RRRRRRRRRqv_1)1 ap_qW1qY__mh  7t_th   7t_v1que_  _ha4Z_X_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 ap_qW1qY__mh  7t_th   7t_v1que_  _ha4Z_X_;u2
R
RRRRRRRRRv1_q1a )_Wqpq_Y1m h_7_t h  t7_t 1uqv_  ehXa_Z__juR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t h  t7_t 1uqv_  ehXa_Z__ju
2;
RRRRRRRRvRR_1q1 _)aqqpWYm1_h7_ t1 _q_vu he aZ_X__XZuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t 1uqv_  ehXa_ZZ_X_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
R
RRRRRRMRC8R

RRRRRHRRVCR58_oC0C$bRR==`pme_Yqh  7t2CRLoRHM:_RlNC##sN0_D$IN#M_F_oC8CM_N$oC8CR
RRRRRRRRRv1_q1a )_Wqpq_Y1m h_7_t q hY7_t uR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t q hY7_t u
2;
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRRRRRqv_1)1 ap_qW1qY__mh  7t_Yqh  7t_1a aX_ uX)_Z:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)qa_pYWq1h_m_t 7 h_qYt 7  _a1 a_X_u)XuZ_2
;
RRRRRRRRR_Rvq 11)qa_pYWq1h_m_t 7 h_qYt 7 q_1v u_ea h__XZuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t q hY7_t 1uqv_  ehXa_Z2_u;R

RRRRRRRRRqv_1)1 ap_qW1qY__mh  7t_Yqh  7t_ u)eq_1v u_ea h__XZuR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_Wqpq_Y1m h_7_t q hY7_t ue) _v1que_  _haXuZ_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRRRRC
M8RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
