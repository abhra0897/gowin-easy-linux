@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)aBpYB  _1Thz B; "
H
`VV8CRpme_QQha1_vtR
RH0MHH
NDRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
HRRMHH0NLDRCMoH
RRRRRHV5lMk_#O	R.<R2CRLo
HMRRRRRPRFDs_Cs_Fs0Q5"DoDCNPDRNCDkRsVFRsbNN0lCCMsRkOl_	I#REEHOR#lk0CRLR0#CRR0FPkNDCsRoCCN0sER0N4MR"
2;RRRRC
M8RMRC8`

HCV8VeRmp]_1q7) _7Bm R

RsbNN0lCChsRB=jRRC5MO#C#N_s$O8FMHF0HM=R=Re`mp)_aQ tt)h_m_1vmaQ_uu; 2
bRRNlsNCs0CR4hBR5=RMCCO#s#N$F_OM08HHRFM=`=Rm_epat)Qt_ )mwh_Qa)1_uuQ 
2;RNRbsCNl0RCshRB.=MR5C#OC#$Ns_MOF8HH0F=MR=mR`eap_)tQt m)_hQ_w)_1ahQmuu; 2
bRRNlsNCs0CRvhz_1Bi_=4RRk5Ml	_O#2-4;R
RbNNslCC0szRhvi_B1R_.=hR5zBv_i41_Rj>R2RR?5vhz_1Bi_-4RRR42:;Rj
R
RsRCorlMk_#O	-j4:9#RRCJJ_kCCk;R
R
HRRMHH0NLDRCMoH
RRRRJ#C_CJkk=CRRk{Ml	_O#'{4L}j};R
RC
M8
NRRD$IN#@R@RF5b#oC8CDRO	L2RCMoH
RRRRRHV5e`mp _)1_ a1hQtq!pR='R4LR42LHCoMR
RRRRR#_CJJkkCC=R<Rk{Ml	_O#'{4L}j};R
RRMRC8R
RRDRC#LCRCMoH
RRRR#RRCJJ_kCCkrlMk_#O	-R49<h=RB?.RR55~|J#C_CJkkMCrkOl_	4#-:2492RR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR&RR&PRCC_M0#kCJCCMOrlMk_#O	-R49:R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRPRCC_M0#kCJCCMOrlMk_#O	-;49
RRRR#RRCJJ_kCCkrvhz_1Bi_j.:9=R<RC5#Jk_JCRkC>4>R2RR&CMPC0C_#JMkCOhCrzBv_i.1_:;j9
RRRR8CM
CRRM
8
`8CMH/VR/eRmp]_1q7) _7Bm `

HCV8VeRmp1_q1a )_
mh
bRRsCFbsR0$q 11)1a_  Tzh_B at)Qt_ )mwh_Qa)1_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRRRFRM0&R55C5#Jk_JCrkCM_klO-	#49:4RC&RP0CM_J#CkOCMCkrMl	_O#:-.jR92|RR
RRRRRRRRR5R~#_CJJkkCCkrMl	_O#:-442922=R!RL4'4R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)a1z T  hB_Qa)t)t __mhvam1_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR#_CJJkkCC9r4R>|-RCCPM#0_CCJkMrOCj
9;RMRC8Fbsb0Cs$


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRFbsb0Cs$1Rq1a )_T1 zB h )_aQ tt)h_m_jhB_4hB_)wQ1 a_ea h__XZuR;
RRRRR5@@bCF#8RoCO2D	
RRRR8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RRRRRH!f#	kMMMFI5CCPM#0_CCJkMrOCM_klO-	#4;92
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 a _1Thz Ba _)tQt m)_hB_h.Q_w)_1a he aZ_X_
u;RRRRR@R@5#bFCC8oR	OD2R
RRRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRRR5R5!#5|CJJ_kCCkrlMk_#O	-44:9R22|f|RHM#k	IMFM|55#_CJJkkCCkrMl	_O#:-442922-R|>R
RRRRR!#fHkMM	F5IMCMPC0C_#JMkCOMCrkOl_	4#-9
2;RRRRCbM8sCFbs
0$
RRRRFbsb0Cs$1Rq1a )_T1 zB h )_aQ tt)h_m_4hB_.hB_A1z1z T _ha he aX1_Z;_u
RRRR@RR@F5b#oC8CDRO	R2
RRRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR!RRfkH#MF	MI5M5^C5#Jk_JCrkCM_klO-	#49:4RC&RP0CM_J#CkOCMCzrhvi_B1:_.j2922R;
RCRRMs8bFsbC0
$
RRRRbbsFC$s0R1q1 _)a1z T  hB_Qa)t)t __mhh_Bjh_mhpaq1_  eh_a1XuZ_;R
RRRRR@b@5F8#CoOCRD
	2RRRRRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRRRR!#fHkMM	F5IM5#^5CJJ_kCCkrlMk_#O	-44:9RR&CMPC0C_#JMkCOhCrzBv_i.1_:Rj9&R
RRRRRRRRRRRRRR{R{5lMk_#O	-{.244'L}{},4j'L}2}22R;
RCRRMs8bFsbC0
$
RRRRbbsFC$s0R1q1 _)a1z T  hB_Qa)t)t __mhh_Bjpaq1_  ehXa_Z__4XuZ_;R
RRRRR@b@5F8#CoOCRD
	2RRRRRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRRRRfkH#MF	MI#M5CJJ_kCCkr249R>|-RR
RRRRR!f5RHM#k	IMFMP5CC_M0#kCJCCMOr2j9RR||CMPC0C_#JMkCOjCr9;R2
RRRR8CMbbsFC$s0
R
RRsRbFsbC0q$R1)1 a _1Thz Ba _)tQt m)_hB_hjq_p1 a_ea h_X4_Z;_u
RRRR@RR@F5b#oC8CDRO	R2
RRRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR5RR!#fHkMM	F5IM#_CJJkkCC9r42|2R-
>RRRRRR5R!#_CJJkkCC9r4RR&&fkH#MF	MICM5P0CM_J#CkOCMC9rj2
2;RRRRCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRh2BjRoLCH:MRRNN_#s#C0C_#JMkCO0C_soHoCFs_MF_l#R0
RRRRRRRRRqq_1)1 a _1Thz Ba _)tQt m)_hm_v1ua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)a1z T  hB_Qa)t)t __mhvam1_Ru2
RRRRRRRRCRRDR#CF_PDCFsss5_0"swH#M0RkOl_	4#-RCCPMR0#FkOOsRC8LRk00$ECRCNsR0MFRDVFDCFI8$RLRC0ER#DN0PRCCRM0H#MRCCJkM"OC2R;
RRRRRCRRMR8
RRRRRHRRVhR5B|4R|BRh.L2RCMoHRN:R_#N#C_s0#kCJCCMO_H0sosoC__FMV#Hs0R
RRRRRRRRRq1_q1a )_T1 zB h )_aQ tt)h_m_)wQ1ua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)a1z T  hB_Qa)t)t __mhw1Q)a2_uRR
RRRRRRRRRCCD#RDFP_sCsF0s_5H"wsR#0CMPC0ORFOCks8kRL00RHRRH#MRF0VDFDF8ICRRL$0RECs0C#RRFV0RECCMPC0H#RMCR#JMkCO2C";R
RRRRRRMRC8`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRH5VRhRBj|h|RB
42RRRRRRRRRCRLoRHM:_RNNC##s#0_CCJkM_OC0osHo_CsFMM_OMj_OV4_H0s#_CCPMG0_xR
RRRRRRRRRR_Rqq 11)1a_  Tzh_B at)Qt_ )mhh_Bhj_Bw4_Qa)1_  ehXa_Z:_u
RRRRRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_jhB_4hB_)wQ1 a_ea h__XZuR2
RRRRRRRRRCRRDR#CF_PDCFsss5_0"swH#C0RP0CMRRHM0REC#kCJCCMORMOF0MNH#RRXFZsR"
2;RRRRRRRRRMRC8R

RRRRRHRRVhR5B
.2RRRRRRRRRCRLoRHM:_RNNC##s#0_CCJkM_OC0osHo_CsFMM_OV._H0s#_CCPMG0_xR
RRRRRRRRRR_Rqq 11)1a_  Tzh_B at)Qt_ )mhh_Bw._Qa)1_  ehXa_Z:_u
RRRRRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_.hB_)wQ1 a_ea h__XZuR2
RRRRRRRRRCRRDR#CF_PDCFsss5_0"swH#C0RP0CMRRHM0REC#kCJCCMORMOF0MNH#RRXFZsR"
2;RRRRRRRRRMRC8R

RRRRRHRRVRR5hRB4|h|RB2.R
RRRRRRRRLRRCMoHRN:R_#N#C_s0#kCJCCMO_H0sosoC__FMM_O4M_O.##kLCCJkMC0_P0CM#x_G
RRRRRRRRRRRRqq_1)1 a _1Thz Ba _)tQt m)_hB_h4B_h.z_1AT1 za h_  eh_a1XuZ_:R
RRRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _1Thz Ba _)tQt m)_hB_h4B_h.z_1AT1 za h_  eh_a1XuZ_2R
RRRRRRRRRRDRC#FCRPCD_sssF_"051#kLCCJkMC0RP0CM#MRHRC0ERJ#CkOCMCFROMH0NMRRXFZsR"
2;RRRRRRRRRMRC8R
RRRRRRRRR
RRRRRRRRRHV5BRhj
R2RRRRRRRRRCRLoRHM:_RNNC##s#0_CCJkM_OC0osHo_CsFMM_OGj_xR
RRRRRRRRRR_Rqq 11)1a_  Tzh_B at)Qt_ )mhh_Bhj_mph_q_1a he aX1_Z:_u
RRRRRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_jhB_hhm_1pqae_  1ha__XZuR2
RRRRRRRRRCRRDR#CF_PDCFsss5_0"swH#M0RkOl_	4#-RCCPMR0#H0MRE#CRCCJkMROCO0FMNRHMXsRFR2Z";R

RRRRRRRRRqRR_1q1 _)a1z T  hB_Qa)t)t __mhh_Bjpaq1_  eh4a___XZuR:
RRRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)1a_  Tzh_B at)Qt_ )mhh_Bpj_q_1a he a__4XuZ_2R
RRRRRRRRRRDRC#FCRPCD_sssF_"05p0N#RCCPMH0RMER0CCR#JMkCOOCRFNM0HRM#XsRFR2Z";R

RRRRRRRRRqRR_1q1 _)a1z T  hB_Qa)t)t __mhh_Bjpaq1_  ehXa_Z__4XuZ_:R
RRRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _1Thz Ba _)tQt m)_hB_hjq_p1 a_ea h__XZ4Z_X_
u2RRRRRRRRRRRRCCD#RDFP_sCsF0s_5H"wsR#0M_klO-	#4PRCC#M0RRHM0REC#kCJCCMORMOF0MNHRFXRs"RZ2R;
RRRRRRRRR8CM
CR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRRHV5jhB2CRLoRHM:_RlNC##s#0_CCJkM_OC0osHo_CsFlM_F
#0RRRRRRRRR_Rvq 11)1a_  Tzh_B at)Qt_ )mvh_m_1auR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_1vma2_u;RR
RRRRRCRRMR8
RRRRRHRRVhR5B|4R|BRh.L2RCMoHRl:R_#N#C_s0#kCJCCMO_H0sosoC__FMV#Hs0R
RRRRRRRRRv1_q1a )_T1 zB h )_aQ tt)h_m_)wQ1ua_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)a1z T  hB_Qa)t)t __mhw1Q)a2_u;RR
RRRRRCRRM
8
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRRHV5jhBRR||h2B4
RRRRRRRRLRRCMoHRl:R_#N#C_s0#kCJCCMO_H0sosoC__FMM_OjM_O4V#Hs0P_CC_M0GRx
RRRRRRRRRvRR_1q1 _)a1z T  hB_Qa)t)t __mhh_Bjh_B4w1Q)ae_  _haXuZ_:R
RRRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a _1Thz Ba _)tQt m)_hB_hjB_h4Q_w)_1a he aZ_X_;u2
RRRRRRRRCRRM
8
RRRRRRRRH5VRh2B.
RRRRRRRRLRRCMoHRl:R_#N#C_s0#kCJCCMO_H0sosoC__FMM_O.V#Hs0P_CC_M0GRx
RRRRRRRRRvRR_1q1 _)a1z T  hB_Qa)t)t __mhh_B.w1Q)ae_  _haXuZ_:R
RRRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a _1Thz Ba _)tQt m)_hB_h.Q_w)_1a he aZ_X_;u2
RRRRRRRRCRRM
8
RRRRRRRRH5VRR4hBRR||hRB.2R
RRRRRRRRRLHCoMRR:l#_N#0Cs_J#CkOCMCs_0HCoosM_F_4MO_.MO_L#k#kCJC_M0CMPC0G#_xR
RRRRRRRRRR_Rvq 11)1a_  Tzh_B at)Qt_ )mhh_Bh4_B1._z A1Thz ae_  1ha__XZuR:
RRRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)1a_  Tzh_B at)Qt_ )mhh_Bh4_B1._z A1Thz ae_  1ha__XZu
2;RRRRRRRRRMRC8R
RRRRRRRRR
RRRRRRRRRHV5BRhj
R2RRRRRRRRRCRLoRHM:_RlNC##s#0_CCJkM_OC0osHo_CsFMM_OGj_xR
RRRRRRRRRR_Rvq 11)1a_  Tzh_B at)Qt_ )mhh_Bhj_mph_q_1a he aX1_Z:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_jhB_hhm_1pqae_  1ha__XZu
2;
RRRRRRRRRRRRqv_1)1 a _1Thz Ba _)tQt m)_hB_hjq_p1 a_ea h_X4_Z:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_jhB_1pqae_  _ha4Z_X_;u2
R
RRRRRRRRRR_Rvq 11)1a_  Tzh_B at)Qt_ )mhh_Bpj_q_1a he aZ_X_X4_Z:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_T1 zB h )_aQ tt)h_m_jhB_1pqae_  _haX4Z___XZu
2;RRRRRRRRRMRC8`
RCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
`

HCV8VeRmpm_Be_ )m
h
RCRoMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RRRRRPOFC#s_CCJkM_OC0osHo:Cs
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	
2RRRRRRRRRRRRRRRRRRRRRR5R5`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRRRRRRRRRRRRRRRRR5h55B|4R|BRh.&2R&PRCC_M0#kCJCCMOrlMk_#O	-249R
||RRRRRRRRRRRRRRRRRRRRRhR5B&jR&#R&CJJ_kCCkr2492
22RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5C"#JMkCO0C_soHoCOsRFsPCC28";R
RRCRRMR8
RCRRM
8
RMRC8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



