-- $Header: //synplicity/map400rc/mappers/xilinx/lib/gen_spartan3/cmp_eq.vhd#1 $
@EH
DLssN$CRHCRC;
Ck#RCHCC03#8F_Do_HO4c4n3DND;C

M00H$JRC_CCDl0CMR
H#RRRRb0Fs5,NjR,LjR,N4R,L4RHD0MRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRR00Fk:kRF00R#8F_Do2HO;M
C8JRC_CCDl0CM;


NEsOHO0C0CksRMCJRRFVCCJ_DCClMH0R##
SHNoMD4R0R#:R0D8_FOoH;

SSlOFbCFMMv0RzYXB_Rp
SFSbs50R
RRRSpSSmRR:FRk0#_08DHFoOR;
RSRSSRBQ:MRHR8#0_oDFH
O;RSRRSQS7RH:RM0R#8F_Do;HO
RRRS1SSRH:RM0R#8F_Do
HOR2SS;C
SMO8RFFlbM0CM;-
S-0N0skHL0#CR$LM_D	NO_GLFRRFVvBzXYR_p:FROlMbFCRM0H0#Rs;kC
oLCHSM
0<4R=NR54MRGFLsR4N2RM58RNGjRMRFsL;j2
RRRRGlk_#HM0RR:vBzXY
_pRRRRRRRRb0FsRblN5=1R>4R0,RR
RRRRRpRRm>R=RFD0k
0,RRRRRRRRB=QR>0RDH
M,RRRRRRRR7=QR>4R''
2;CRM8C;JM
D

HNLssH$RC;CCR#
kCCRHC#C30D8_FOoH_n44cD3ND
;
CHM00C$RJD_CCMlC0M_FC0LHR
H#RRRRb0Fs5,NjR,LjRHD0MRR:H#MR0D8_FOoH;R
RRRRRRRRRRDRR00Fk:kRF00R#8F_Do2HO;M
C8JRC_CCDl0CM_CFML;H0
N

sHOE00COkRsCCRJMFCVRJD_CCMlC0M_FC0LHR
H#So#HMRND0:4RR8#0_oDFH
O;SO
SFFlbM0CMRXvzBpY_
SRSb0FsRR5
RSRSSRpm:kRF00R#8F_Do;HO
RRRSBSSQRR:H#MR0D8_FOoH;R
RRSSS7:QRRRHM#_08DHFoOR;
RSRSS:1RRRHM#_08DHFoOS
RS
2;S8CMRlOFbCFMM
0;SN--0H0sLCk0RM#$_NLDOL	_FFGRVzRvX_BYpRR:ObFlFMMC0#RHRk0sCL;
CMoH
4S0RR<=5RNjGsMFR2Lj;R
RRkRlGM_H#:0RRXvzBpY_
RRRRRRRRsbF0NRlbR51=0>R4
,RRRRRRRRRp=mR>0RDF,k0
RRRRRRRRRBQ=D>R0,HM
RRRRRRRRR7Q='>R4;'2
8CMRMCJ;



LDHs$NsRCHCC
;RkR#CHCCC38#0_oDFH4O_43ncN;DD
M
C0$H0RuBv_R THR#
RoRRCsMCHIO5HE80RH:RMo0CC:sR=;42
RRRRsbF0:5qRRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRR:RARRHM#_08DHFoOC_POs0F58IH0-ER4FR8IFM0R;j2
RRRRRRRRTR RF:Rk#0R0D8_FOoH2C;
MB8Rv u_T
;

ONsECH0Os0kCCRODDD_CDPCRRFVB_vu HTR#V

k0MOHRFMVOkM_sCsFCs5JH_I8R0E:MRH0CCoss2RCs0kM0R#soHMR
H#LHCoMR
RH5VR5_CJI0H8E=R>R24.R8NMRJ5C_8IH0<ER=cRn202RE
CMRRRRskC0s"M5"
2;RDRC#RC
RsRRCs0kMC5"sssF"
2;RMRC8VRH;M
C8kRVMCO_sssF;0
N0LsHkR0CoCCMsFN0sC_sb0FsR#:R0MsHoN;
0H0sLCk0RMoCC0sNFss_CsbF0VRFRDOCDC_DPRCD:sRNO0EHCkO0sHCR#kRVMCO_sssF58IH0;E2
O
SF0M#NRM0Hs0CNF0HMRR:HCM0oRCs:5=RI0H8E.2/;O
SF0M#NRM0sNClHCM8sRR:HCM0oRCs:5=RI0H8El2RF.8R;R
RRHR#oDMNR08NNl_0bRR:#_08DHFoOC_POs0FRH5I8R0E-RR48MFI0jFR2S;
#MHoNhDR :TRR8#0_oDFH
O;SR
RRFROlMbFCRM0CCJ_DCClMH0R#R
RRRRRRFRbsN05jL,RjN,R4L,R4D,R0:HMRRHM#_08DHFoOR;
RRRRRRRRRRRRRRRRDk0F0RR:FRk0#_08DHFoO
2;RRRRCRM8ObFlFMMC0
;
SlOFbCFMMC0RJD_CCMlC0M_FC0LHR
H#RRRRRRRRb0Fs5,NjR,LjRHD0MH:RM0R#8F_Do;HO
RRRRRRRRRRRRRRRR0RDFRk0:kRF00R#8F_Do2HO;R
RRMRC8FROlMbFC;M0
oLCHSM
z:jRR5HVR8IH0>ERRR42oCCMsCN0
CSLo
HMRRRRzRj4:JRC_CCDl0CM
RRRRRRRRRRRRRRRRsbF0NRlbS5
SNSSj>R=Rjq52
,RRRRRRRRRRRRRRRRRL=jR>5RAj
2,SSSSN=4R>5Rq4R2,
RRRRRRRRRRRRRRRRRL4=A>R5,42
RRRRRRRRRRRRRRRRHD0M>R=R''j,R
RRRRRRRRRRRRRR0RDFRk0=8>RN_0N05lbj;22
MSC8CRoMNCs0
C;
RRRRRRRRz
S4RR:HRV5I0H8ERR=4o2RCsMCN
0CSoLCHSM
STh RR<=q25jRFGMs5RAj
2;S8CMRMoCC0sNC
;
RRRRz:.RRsVFR0LH_8HMCHGRMRR405FRHs0CNF0HMRR-4R2RoCCMsCN0
RRRRRRRRoLCHRM
RRRRRRRRRzRR.:4RR_CJClDCC
M0RRRRRRRRRRRRRRRRb0FsRblN5S
SSjSNRR=>q*5.L_H0HCM8GR2,
RRRRRRRRRRRRRRRRRLj=A>R5L.*HH0_MG8C2S,
SNSS4>R=R.q5*0LH_8HMC+GRR,42RR
RRRRRRRRRRRRRR4RLRR=>A*5.L_H0HCM8GRR+4
2,RRRRRRRRRRRRRRRRDM0HRR=>8NN0_b0l50LH_8HMC-GRR,42
RRRRRRRRRRRRRRRRFD0k=0R>NR800N_lLb5HH0_MG8C2
2;RRRRRRRRCRM8oCCMsCN0;S

z:dRR5HVRlsCN8HMC=sRRN4RMI8RHE80R4>R2CRoMNCs0SC
LHCoMS
SzRd4:JRC_CCDl0CM_CFML
H0SbSSFRs0l5Nb
SSSSRNj=q>R58IH0-ER4
2,SSSSL=jR>5RAI0H8ERR-4
2,SSSSDM0HR8=>N_0N05lbHs0CNF0HMRR-4
2,SSSSDk0F0>R=RTh 2S;
CRM8oCCMsCN0;R

RRRRR
RRSRzc:VRH5lsCN8HMC=sRRNjRMI8RHE80RRR>4o2RCsMCN
0CSoLCHRM
RSRRhR T<8=RN_0N05lbHs0CNF0HMRR-4R2;
C
SMo8RCsMCN;0C
SS
zR6: <TR=FRM0 5hT
2;
8CMRCRODDD_CDPC;



