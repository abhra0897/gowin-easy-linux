`ifndef ATCWDT200_CONST_VH
`define ATCWDT200_CONST_VH

`define ATCWDT200_PRODUCT_ID		32'h03002004

`endif

