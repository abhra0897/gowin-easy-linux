@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Ta_z1Q Ba h_q1aa; "
R
R`OHMDCk8R0"#8P_FDN_0#E	3"


`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/eRmph_QQva_1
t
`8HVCmVReqp_1)1 ah_m
H
`VV8CRpme_7 h__mw1zQvpQqamRh
RbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aau _;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRfR5sCF#5e`mph_ 7w_m_v1QzapqQ2mhR
||RRRRRFfs##C5NDlbCP_CC2M02-R|>#R50CN0_bCGs=R=RCOEOP	_NCDk2R;
RCRRMs8bFsbC0
$
RHR`VV8CRpme_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRRR/R/7MFRFH0EMRo
R`RRCCD#
RRRRbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aaX _Zh_m_1 m_
u;RRRRR@R@5#bFCC8oR	OD2R
RRRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRRR5R5!H5f#	kMMMFI5b5fN5#0`pme_7 h__mw1zQvpQqam2h22&2R&5R!5Nfb#`05m_ep _h7m1w_QpvzqmaQh222RR
RRRRRR&R&Rf!5HM#k	IMFMm5`e p_hm7_wQ_1vqzpahQm2R22|R|
RRRRR!R55#fHkMM	F5IM5Nfb#`05m_ep _h7m1w_QpvzqmaQh2222&R&Rf55b0N#5e`mph_ 7w_m_v1QzapqQ2mh2R22|R|
RRRRR5R5fkH#MF	MI5M5f#bN0m5`e p_hm7_wQ_1vqzpahQm2222RR&&!H5f#	kMMMFI5e`mph_ 7w_m_v1QzapqQ2mh2R
RRRRRR&RR&5R!`pme_7 h__mw1zQvpQqamRh22
2;RRRRRMRC8Fbsb0Cs$R

RRRRRFbsb0Cs$1Rq1a )_QTz  1Bh1a_a qa__XZm1h_a qa_u X);_u
RRRR@RR@F5b#oC8CDRO	R2
RRRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR5RRf#sFCm5`e p_hm7_wQ_1vqzpahQm2|R|
RRRRRRRRRRRRsRfF5#C#bNlDCC_P0CM2|2R-5>R!H5f#	kMMMFI5N#00CC_G2bs2
2;RRRRRMRC8Fbsb0Cs$R

RRRRRFbsb0Cs$1Rq1a )_QTz  1Bh1a_a qa__XZmBh_]i B_peqzu _;R
RRRRR@b@5F8#CoOCRD
	2RRRRRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRRRR5Ffs#`C5m_ep _h7m1w_QpvzqmaQh|2R|R
RRRRRRFfs##C5NDlbCP_CC2M02-R|>!R55#fHkMM	F5IMOOEC	N_PD2kC2
2;RRRRRMRC8Fbsb0Cs$R
RRCR`MV8HRm//eQp_vQupB_QaX B]Bmi_wRw
RM`C8RHV/e/mpB_X]i B_wmw
D`C#RC
RbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aau _;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRsRfF5#C#bNlDCC_P0CM2-R|>#R50CN0_bCGs=R=RCOEOP	_NCDk2R;
RCRRMs8bFsbC0
$
RHR`VV8CRpme_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRRR/R/7MFRFH0EMRo
R`RRCCD#
RRRRbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aaX _Zh_m_q1aa  _X_u)uR;
RRRRR5@@bCF#8RoCO2D	
RRRR8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RRRRRFfs##C5NDlbCP_CC2M0R>|-R55!fkH#MF	MI#M50CN0_bCGs222;R
RRRRRCbM8sCFbs
0$
RRRRbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aaX _Zh_m_ B]Bei_q pz_
u;RRRRR@R@5#bFCC8oR	OD2R
RRRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRRRsRfF5#C#bNlDCC_P0CM2-R|>!R55#fHkMM	F5IMOOEC	N_PD2kC2
2;RRRRRMRC8Fbsb0Cs$R
RRM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mw`
RCHM8V/R/m_epX B]Bmi_w`w
CHM8V/R/Rpme_7 h__mw1zQvpQqam
h
`8HVCmVReXp_BB] iw_mwR
RR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RbRRsCFbsR0$q 11)Ta_z1Q Ba h_q1aaX _Zh_m_v1qu_p  he a;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR!555#fHkMM	F5IM5Nfb##05NDlbCP_CC2M02R22&!&R5b5fN5#0#bNlDCC_P0CM2R22
RRRR&RR&5R!fkH#MF	MI#M5NDlbCP_CC2M02|2R|R
RR5RR!H5f#	kMMMFI5b5fN5#0#bNlDCC_P0CM2222RR&&5b5fN5#0#bNlDCC_P0CM2222R
||RRRRRf55HM#k	IMFMf55b0N#5l#Nb_DCCMPC02222&R&Rf!5HM#k	IMFMN5#lCbD_CCPM202
RRRRRRR&!&R5l#Nb_DCCMPC022R2R;
RCRRMs8bFsbC0R$
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)aT zQ1hB aa_1q_a uN:R#s#C0sRbFsbC05$Rq 11)Ta_z1Q Ba h_q1aau _2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05100NCGRCb#sC#MHFRRH#MRF0CNJkDFR0RCOEOP	_NCDkRHIED#CRNDlbCPRCCRM0HN#R#s#C0"C82
;
RRRR`8HVCmVReXp_BB] iw_mwR
RRRRRR/R/7MFRFH0EMRo
R`RRCCD#
RRRR`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RRRRRR/R/7MFRFH0EMRo
RRRRRD`C#RC
RRRRRqRR_1q1 _)aT zQ1hB aa_1q_a XmZ_ha_1q_a  )Xu_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)aT zQ1hB aa_1q_a XmZ_ha_1q_a  )Xu_
u2RRRRRRRRCCD#RDFP_sCsF0s_50"#N_0CCsGbRMOF0MNH#RRXFZsR"
2;
RRRRRRRRqq_1)1 az_TQB 1 _ha1aaq Z_X__mhBB] iq_ep_z uR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)Ta_z1Q Ba h_q1aaX _Zh_m_ B]Bei_q pz_
u2RRRRRRRRCCD#RDFP_sCsF0s_5E"OC_O	PkNDCFROMH0NMX#RRRFsZ;"2
R
RRRRRR_Rqq 11)Ta_z1Q Ba h_q1aaX _Zh_m_v1qu_p  he a:_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_QTz  1Bh1a_a qa__XZm1h_qpvu e_  _hauR2
RRRRRCRRDR#CF_PDCFsss5_0"l#Nb_DCCMPC0FROMH0NMX#RRRFsZ;"2
R
RRRRRRHR`VV8CRpme_7 h__mw1zQvpQqamRh
RRRRRRRRRqq_1)1 az_TQB 1 _ha1aaq Z_X__mh _m1uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_QTz  1Bh1a_a qa__XZm h_mu1_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5m"`e p_hm7_wQ_1vqzpahQmRMOF0MNH#RRXFZsR"
2;RRRRRRRR`8CMH/VR/pme_7 h__mw1zQvpQqam
h
RRRRRCR`MV8HRm//eQp_vQupB_QaX B]Bmi_wRw
R`RRCHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 az_TQB 1 _ha1aaq :_uR#N#kRlCbbsFC$s0R15q1a )_QTz  1Bh1a_a qa_;u2
R
RRHR`VV8CRpme_]XB _Bim
wwRRRRRRRR/F/7R0MFEoHM
RRRRD`C#RC
RRRRRV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRRRRRR/F/7R0MFEoHM
RRRR`RRCCD#
RRRRRRRRqv_1)1 az_TQB 1 _ha1aaq Z_X__mh1aaq X_ uu)_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 az_TQB 1 _ha1aaq Z_X__mh1aaq X_ uu)_2
;
RRRRRRRRv1_q1a )_QTz  1Bh1a_a qa__XZmBh_]i B_peqzu _:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 az_TQB 1 _ha1aaq Z_X__mhBB] iq_ep_z u
2;
RRRRRRRRqv_1)1 az_TQB 1 _ha1aaq Z_X__mh1uqvp  _ea h_
u:RRRRRRRRNk##lbCRsCFbsR0$51q1 _)aT zQ1hB aa_1q_a XmZ_hq_1v up_  ehua_2
;
RRRRRRRR`8HVCmVRe p_hm7_wQ_1vqzpahQm
RRRRRRRRvRR_1q1 _)aT zQ1hB aa_1q_a XmZ_hm_ 1:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)Ta_z1Q Ba h_q1aaX _Zh_m_1 m_;u2
RRRRRRRRM`C8RHV/e/mph_ 7w_m_v1QzapqQ
mh
RRRR`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
wwRRRR`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m




