`ifndef ATCPIT100_CFG_VH
`define ATCPIT100_CFG_VH
`include "ae250_config.vh"
`include "ae250_const.vh"
//-------------------------------------------------
// Number of PIT Channels
//-------------------------------------------------
//`define ATCPIT100_NUM_CHANNEL_1
//`define ATCPIT100_NUM_CHANNEL_2
//`define ATCPIT100_NUM_CHANNEL_3
//`define ATCPIT100_NUM_CHANNEL_4

`endif // ATCPIT100_CFG_VH
