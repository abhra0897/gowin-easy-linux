@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Qa_vQupBQqam;h"
R
R`OHMDCk8R0"#8P_FDN_0#E	3"


`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vt`

HCV8VeRmp1_q1a )_
mh
bRRsCFbsR0$q 11)Qa_vQupBQqamuh_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RNCM0OCC8MC0_GRbs|R->O#FMCCJkMC0_G;bs
CRRMs8bFsbC0
$

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RbbsFC$s0R1q1 _)aQpvuQaBqQ_mhXmZ_hh_qaX_ u;_u
@RR@bR5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5HM#k	IMFMM5N0CCO80CM_bCGs222;R
RCbM8sCFbsR0$
R
RbbsFC$s0R1q1 _)aQpvuQaBqQ_mhXmZ_hm_BhX_ u;_u
@RR@bR5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RNCM0OCC8MC0_GRbs|R->5f!5HM#k	IMFMF5OMJ#Ck0CM_bCGs222;R
RCbM8sCFbsR0$
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
oRRCsMCN
0C
RRRR#ONCbR5sCFbs_0$0C$b2R
RRRRR`pme_1q1 R)a:CRLoRHM:PRFD#_N#0Cs
RRRRRRRRqq_1)1 av_QuBpQqmaQh:_uR#N#CRs0bbsFC$s0R15q1a )_uQvpqQBahQm_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RDFP_sCsF0s_5M"q0CCO80CMRC8F#FRM0NREPOCRFCM#JMkC0;"2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRqRR_1q1 _)aQpvuQaBqQ_mhXmZ_hh_qaX_ u:_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_uQvpqQBahQm__XZmqh_h a_Xuu_2R
RRRRRRDRC#FCRPCD_sssF_"05NCM0OCC8MC0_GRbsO0FMN#HMRFXRs"RZ2R;
RRRRR
RRRRRRRRRRq1_q1a )_uQvpqQBahQm__XZmBh_m h_Xuu_:R
RRRRRR#RN#0CsRFbsb0Cs$qR51)1 av_QuBpQqmaQhZ_X__mhB_mh _XuuR2
RRRRRCRRDR#CF_PDCFsss5_0"MOF#kCJC_M0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRv1_q1a )_uQvpqQBahQm_Ru:Nk##lbCRsCFbsR0$51q1 _)aQpvuQaBqQ_mhu
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rvq 11)Qa_vQupBQqamXh_Zh_m_aqh_u X_
u:RRRRRRRRNk##lbCRsCFbsR0$51q1 _)aQpvuQaBqQ_mhXmZ_hh_qaX_ u2_u;R
RRRRRRRR
RRRRRvRR_1q1 _)aQpvuQaBqQ_mhXmZ_hm_BhX_ u:_u
RRRRRRRR#N#kRlCbbsFC$s0R15q1a )_uQvpqQBahQm__XZmBh_m h_Xuu_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epQmth): RRoLCH:MRRDFP_MHoF
sCRRRRRRRR/8/RFFRM0MEHoR
RRRRRC
M8RR
RRRRR8NCVkRD0RRRR:MRHHN0HDPRFDs_Cs_Fs0"5"2R;
RCRRMN8O#
C
RMRC8MoCC0sNC`

CHM8V/R/Rpme_1q1 _)am
h
`8HVCmVReBp_m)e _
mh
oRRCsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_CsNCM0OCC8M
0:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRNCM0OCC8MC0_G2bsRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"0NMC8OCCRM0OCFPs"C82
;
RRRRR8CM
RRRR8CM
R
RCoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
