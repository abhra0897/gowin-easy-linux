
@ER--=========m==F=FF=========================================FmFF========-
-RR=RB$FbsEHo0BR52jR.4.c-jR4gtHFIMCR1lFHOMO8k0RFsaECOMFFDoB$RFp3,0
83-=-RRRRRRRRRRRRRRRRRRRRRRDqDRosHER0#sCC#s8PC3-
-R====================================================================-=
--
-R_R_RRRRR_R_RRRRR_R_
R--R\\RRRRR/\RRRRRR/RR/RwRrHRDCMCNlR9RRRHbsl$_#ME3P8-
-R\RRRR\R/\R/RR\R/RR/RrRR7OC#s0HbHRFM9WRtdRqaep]7RMVkOF0HMRND#0$MEHC##HRDLssN$-
-RRRR\/R\RR/R\/R\RR/RRrRRaCHl#l0NbRRR9CRW8NRvsROEn4R4::jjd.jRj
4g-R-RR\RRRRR/R\RRRRR/RRRRRCrPsF#HMRRRRRR94
34-R-RRRRR\R/RRRRR\R/RRRRRR-
-
R--=========m==F=FF=========================================FmFF========


-------------------------b--NNO	ooCRDNFLD----------------------------
--
ApQ)Yq)RCHCC
;RzR1 HCCC38#0_oDFH4O_43ncN;DDR#
kC RQ 1 3ap7_mBtQ_Qq)aq]3p
p;kR#CQ   371a_tpmQzB_ht1Qh3 7q;pp
q
uBtiq FROlMbFC#M0RRQ1
RRRNs00H0LkC$R#MD_LN_O	L:FGRFLFDMCNRR;
R0RN0LsHkR0C#_$MLODN	F_LGVRFRlBFbCFMMR0#:NRbOo	NC#RHRk0sCR;
R0RN0LsHkR0CLODN	F_LGN_b8H_bM#:R0MsHoR;
R0RN0LsHkR0C#_$MMsFbkRMC:FRLFNDCMR;
R0RN0LsHkR0CGlO_NRb:#H0sM
o;RNRR0H0sLCk0R_GOlRNbFBVRFFlbM0CM#RR:b	NONRoCH"#RD"k0;
RS-----------------------------1-t)---------------------------------------
m
Bvhum RhatR1)
RRRR)uma
R5RRRRRRRRtQ1)RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFtVR1:)RRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkC$R#MF_MbMskCVRFR)t1RB:RFFlbM0CMRRH#0Csk;-

-------------------------apz4----------------------------
--Bumvmhh azRpa
4RRRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"Rj"2R;
RuRRmR)a5R
RRRRRRRRw:kRF00R#8F_Do;HO
RRRRRRRRRQj:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRapz4RR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0R_GOlRNbFpVRzRa4:FROlMbFCRM0H"#RD"k0;

S-------------------------z-pa-.R----------------------------
vBmu mhhpaRzRa.
RRRRht  B)QR
5RRRRRRRRRQahQRL:RHP0_CFO0s=R:RjX""RR
R2RR;R
RRmRu)5aR
RRRSRRRR:wRR0FkR8#0_oDFH
O;RSRRRRRRQ:jRRRHM#_08DHFoOR;
RRRSRQRR4RR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVp.zaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRa.:FROlMbFCRM0H"#RD"k0;-

-------------------------apzd----------------------------
--Bumvmhh azRpa
dRRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0C_POs0FRR:=Xj"j"RR
R2RR;R
RRmRu)5aR
RRRSRRRR:wRR0FkR8#0_oDFH
O;RSRRRRRRQ:jRRRHM#_08DHFoOR;
RRRSRQRR4RR:H#MR0D8_FOoH;R
RRRSRR.RQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:dRRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapzdRR:ObFlFMMC0#RHRk"D0
";
------------------------p--zRac-----------------------------m
Bvhum RhapczaRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:L_H0P0COF:sR="RXjjjj"RR
R2RR;R
RRmRu)5aR
RRRSRRRR:wRR0FkR8#0_oDFH
O;RSRRRRRRQ:jRRRHM#_08DHFoOR;
RRRSRQRR4RR:H#MR0D8_FOoH;R
RRRSRR.RQRH:RM0R#8F_Do;HO
RRRSRRRRRQd:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRapzcRR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVpczaRO:RFFlbM0CMRRH#"0Dk"R;
R
RR-------------------------z-pa-6R----------------------------
vBmu mhhpaRzRa6
RRRRht  B)QR
5RRRRRRRRRQahQRL:RHP0_CFO0s=R:RjX"jjjjj"jjRR
RR;R2
RRRR)uma
R5RSRRRRRRwRR:FRk0#_08DHFoOR;
RRRSRQRRjRR:H#MR0D8_FOoH;R
RRRSRR4RQRH:RM0R#8F_Do;HO
RRRSRRRRRQ.:MRHR8#0_oDFH
O;RSRRRRRRQ:dRRRHM#_08DHFoOR;
RRRSRQRRcRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRa6:FRBlMbFCRM0H0#Rs;kC
0SN0LsHkR0CGlO_NFbRVzRpa:6RRlOFbCFMMH0R#DR"k;0"
RRRR-
-------------------------pnzaR----------------------------B-
mmvuha hRapznRR
RtRR )h Q5BRRR
RRRRRRhRQQ:aRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjj
"RRRRR2R;
RuRRmR)a5R
RRRSRRRRw:kRF00R#8F_Do;HO
RRRSRRRRRQj:MRHR8#0_oDFH
O;RSRRRRRRQ:4RRRHM#_08DHFoOR;
RRRSRQRR.RR:H#MR0D8_FOoH;R
RRRSRRdRQRH:RM0R#8F_Do;HO
RRRSRRRRRQc:MRHR8#0_oDFH
O;RSRRRRRRQ:6RRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVpnzaRB:RFFlbM0CMRRH#0Csk;N
S0H0sLCk0R_GOlRNbFpVRzRan:FROlMbFCRM0H"#RD"k0;-

-------------------------apz(-R--------------------------
--
vBmu mhhpaRzRa(
RRRRht  B)QR
5RRRRRRRRRQahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRR
RR;R2
RRRR)uma
R5RSRRRRRRwRR:FRk0#_08DHFoOR;
RRRSRQRRjRR:H#MR0D8_FOoH;R
RRRSRR4RQRH:RM0R#8F_Do;HO
RRRSRRRRRQ.:MRHR8#0_oDFH
O;RSRRRRRRQ:dRRRHM#_08DHFoOR;
RRRSRQRRcRR:H#MR0D8_FOoH;R
RRQRS6RR:H#MR0D8_FOoH;R
RRRSRRnRQRH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:(RRlBFbCFMMH0R#sR0k
C;S0N0skHL0GCRON_lbVRFRapz(RR:ObFlFMMC0#RHRk"D0
";
------------------------p--zRaU-----------------------------m
Bvhum RhapUzaRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR
R2RR;R
RRmRu)5aR
RRRSRRRR:wRR0FkR8#0_oDFH
O;RSRRRRRRQ:jRRRHM#_08DHFoOR;
RRRSRQRR4RR:H#MR0D8_FOoH;R
RRRSRR.RQRH:RM0R#8F_Do;HO
RRRSRRRRRQd:MRHR8#0_oDFH
O;RSRRRRRRQ:cRRRHM#_08DHFoOR;
RRRSRQRR6RR:H#MR0D8_FOoH;R
RRRSRRnRQRH:RM0R#8F_Do;HO
RRRSRRRRRQ(:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRapzURR:BbFlFMMC0#RHRk0sCS;
Ns00H0LkCORG_blNRRFVpUzaRO:RFFlbM0CMRRH#"0Dk"
;
-------------------------z-vX-.-----------------------------
vBmu mhhvaRzRX.
RRRR)uma
R5SRRRRRQj:MRHR8#0_oDFH
O;SRRRRRQ4:MRHR8#0_oDFH
O;SRRRRR1j:MRHR8#0_oDFH
O;SRRRR:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.RR:BbFlFMMC0#RHRk0sC
;
-------------------------z-vXp._z-a6-----------------------------m
Bvhum Rhav.zX_apz6RR
RuRRmR)a5R
SRQRRjRR:H#MR0D8_FOoH;R
SRQRR4RR:H#MR0D8_FOoH;R
SR1RRjRR:H#MR0D8_FOoH;R
SRmRRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.p6zaRB:RFFlbM0CMRRH#0Csk;-

-------------------------Xvz.z_pa-n-----------------------------
vBmu mhhvaRz_X.pnzaRR
RRmRu)5aR
RSRRjRQRH:RM0R#8F_Do;HO
RSRR4RQRH:RM0R#8F_Do;HO
RSRRjR1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRan:FRBlMbFCRM0H0#Rs;kC
-
-------------------------v.zX_apz(----------------------------
--Bumvmhh azRvXp._zRa(
RRRR)uma
R5SRRRRRQj:MRHR8#0_oDFH
O;SRRRRRQ4:MRHR8#0_oDFH
O;SRRRRR1j:MRHR8#0_oDFH
O;SRRRR:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_pa:(RRlBFbCFMMH0R#sR0k
C;
------------------------v--z_X.pUza-----------------------------B-
mmvuha hRXvz.z_pa
URRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRR1:jRRRHM#_08DHFoOS;
RRRRmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apzURR:BbFlFMMC0#RHRk0sC
;
-------------------------z-vXv._z-XU-----------------------------m
Bvhum Rhav.zX_XvzURR
RuRRmR)a5R
SRQRRjRR:H#MR0D8_FOoH;R
SRQRR4RR:H#MR0D8_FOoH;R
SR1RRjRR:H#MR0D8_FOoH;R
SRmRRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRz_X.vUzXRB:RFFlbM0CMRRH#0Csk;-

-------------------------Xvz.z_vX-4n-----------------------------m
Bvhum Rhav.zX_Xvz4
nRRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRR1:jRRRHM#_08DHFoOS;
RRRRmRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_Xvz4:nRRlBFbCFMMH0R#sR0k
C;
------------------------v--z_X.vdzX.----------------------------
--Bumvmhh azRvXv._z.XdRR
RRmRu)5aR
RSRRjRQRH:RM0R#8F_Do;HO
RSRR4RQRH:RM0R#8F_Do;HO
RSRRjR1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXv._z.XdRB:RFFlbM0CMRRH#0Csk;R
RR-R
-------------------------Xvzc----------------------------
--Bumvmhh azRvX
cRRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRRQ:.RRRHM#_08DHFoO
;RSRRRRRQd:MRHR8#0_oDFH
O;SRRRRR1j:MRHR8#0_oDFH
O;SRRRRR14:MRHR8#0_oDFH
O;SRRRR:mRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzcRR:BbFlFMMC0#RHRk0sC
;
-------------------------z-vX-U-----------------------------
vBmu mhhvaRzRXU
RRRR)uma
R5SRRRRRQj:MRHR8#0_oDFH
O;SRRRRRQ4:MRHR8#0_oDFH
O;SRRRRRQ.:MRHR8#0_oDFHRO;
RSRRdRQRH:RM0R#8F_Do;HO
RSRRcRQRH:RM0R#8F_Do;HO
RSRR6RQRH:RM0R#8F_Do;HO
RSRRnRQRH:RM0R#8F_Do;HO
RSRR(RQRH:RM0R#8F_Do;HO
RSRRjR1RH:RM0R#8F_Do;HO
RSRR4R1RH:RM0R#8F_Do;HO
RSRR.R1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvX:URRlBFbCFMMH0R#sR0k
C;
------------------------v--znX4-----------------------------m
Bvhum Rhav4zXn
RRRRRRuam)RS5
RRRRQ:jRRRHM#_08DHFoOS;
RRRRQ:4RRRHM#_08DHFoOS;
RRRRQ:.RRRHM#_08DHFoO
;RSRRRRRQd:MRHR8#0_oDFH
O;SRRRRRQc:MRHR8#0_oDFH
O;SRRRRRQ6:MRHR8#0_oDFH
O;SRRRRRQn:MRHR8#0_oDFH
O;SRRRRRQ(:MRHR8#0_oDFH
O;SRRRRRQU:MRHR8#0_oDFH
O;SRRRRRQg:MRHR8#0_oDFH
O;SRRRRjQ4RH:RM0R#8F_Do;HO
RSRR4RQ4RR:H#MR0D8_FOoH;R
SRQRR4:.RRRHM#_08DHFoOS;
RRRRQR4d:MRHR8#0_oDFH
O;SRRRRcQ4RH:RM0R#8F_Do;HO
RSRR4RQ6RR:H#MR0D8_FOoH;R
SR1RRjRR:H#MR0D8_FOoH;R
SR1RR4RR:H#MR0D8_FOoH;R
SR1RR.RR:H#MR0D8_FOoH;R
SR1RRdRR:H#MR0D8_FOoH;R
SRmRRRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFvVRznX4RB:RFFlbM0CMRRH#0Csk;-

-------------------------Xvzd-.--------------------------
--Bumvmhh azRvXRd.RR
RRmRu)5aR
RSRRjRQRH:RM0R#8F_Do;HO
RSRR4RQRH:RM0R#8F_Do;HO
RSRR.RQRH:RM0R#8F_Do;HORR
SRQRRdRR:H#MR0D8_FOoH;R
SRQRRcRR:H#MR0D8_FOoH;R
SRQRR6RR:H#MR0D8_FOoH;R
SRQRRnRR:H#MR0D8_FOoH;R
SRQRR(RR:H#MR0D8_FOoH;R
SRQRRURR:H#MR0D8_FOoH;R
SRQRRgRR:H#MR0D8_FOoH;R
SRQRR4:jRRRHM#_08DHFoOS;
RRRRQR44:MRHR8#0_oDFH
O;SRRRR.Q4RH:RM0R#8F_Do;HO
RSRR4RQdRR:H#MR0D8_FOoH;R
SRQRR4:cRRRHM#_08DHFoOS;
RRRRQR46:MRHR8#0_oDFH
O;SRRRRnQ4RH:RM0R#8F_Do;HO
RSRR4RQ(RR:H#MR0D8_FOoH;R
SRQRR4:URRRHM#_08DHFoOS;
RRRRQR4g:MRHR8#0_oDFH
O;SRRRRjQ.RH:RM0R#8F_Do;HO
RSRR.RQ4RR:H#MR0D8_FOoH;R
SRQRR.:.RRRHM#_08DHFoOS;
RRRRQ:.dRMRHR8#0_oDFH
O;SRRRRcQ.RH:RM0R#8F_Do;HO
RSRR.RQ6RR:H#MR0D8_FOoH;R
SRQRR.:nRRRHM#_08DHFoOS;
RRRRQR.(:MRHR8#0_oDFH
O;SRRRRUQ.RH:RM0R#8F_Do;HO
RSRR.RQgRR:H#MR0D8_FOoH;R
SRQRRd:jRRRHM#_08DHFoOS;
RRRRQRd4:MRHR8#0_oDFHRO;
RSRRjR1RH:RM0R#8F_Do;HO
RSRR4R1RH:RM0R#8F_Do;HO
RSRR.R1RH:RM0R#8F_Do;HO
RSRRdR1RH:RM0R#8F_Do;HO
RSRRcR1RH:RM0R#8F_Do;HO
RSRRRRm:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXRd.:FRBlMbFCRM0H0#Rs;kC
-
-------------------------q-pz-----------------------------B-
mmvuha hRzqpRR
RR RthQ )BRR5RR
SRqRRpvz_mR7 :hRQa  t)=R:R
j;RRRRRRRRqR77:hRQa  t)=R:R;jR
RRRRRRRSA1zRQ:Rhta  :)R=RR4;R
RRRRRR7Rq7A1zRQ:Rhta  :)R=RR.;R
RRRRRR ShRQ:Rhta  :)R=RRd;R
RRRRRR StRQ:Rhta  :)R=RRc;R
SRpRR RR:Q hatR ):6=R;R
RRRRRRzSBuRR:Q hatR ):n=RRR;
RRRRRBRR7:hRRaQh )t RR:=(
R;RRRRRRRRBBzu7:hRRaQh )t RR:=US;
RRRRvazpRQ:Rhta  :)R=
RgRRRR2
;SRRRRuam)RS5
RRRR1Rzv:zRma0R#8F_Do;HO
RSRRmRBz:aRRamzR8#0_oDFHSO;
RSRRjRQRQ:Rh0R#8F_Do;HO
RSRR4RQ:hRQR8#0_oDFH
O;SRRRR:QdRRQh#_08DHFoOS;
RRRRB:QhRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRzqpRB:RFFlbM0CMRRH#0Csk;-

-------------------------7--w-wR-----------------------------m
Bvhum Rha7Rww
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''R
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HOSR
SRBRRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wRB:RFFlbM0CMRRH#0Csk;-

-------------------------w-7w- R--------------------------------
vBmu mhh7aRwRw 
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRBRR RR:Q#hR0D8_FOoH;SS
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w: RRlBFbCFMMH0R#sR0k
C;
------------------------w-7w-1R--------------------------------
vBmu mhh7aRwRw1
RRRRht  B)QR
5RRRRRRRRRQahQ:HRL0=R:R''4RR
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HO
RSRR R1aRR:Q#hR0D8_FOoH;SS
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:1RRlBFbCFMMH0R#sR0k
C;
----------------------------w7w1- -------------------------------------
vBmu mhh7aRw w1RR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=R4R'
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;R
SR7RRRQ:Rh0R#8F_Do;HO
RSRR R1aRR:Q#hR0D8_FOoH;R
SRBRR Q:Rh0R#8F_Do;HO
RSRRpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV71ww RR:BbFlFMMC0#RHRk0sC
;
------------------------7)wwR--------------------------------
--Bumvmhh awR7w
)RRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''j
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFH
O;SRRRR:7RRRQh#_08DHFoOS;
RRRR)  1aRR:Q#hR0D8_FOoH;R
SRBRRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w)RR:BbFlFMMC0#RHRk0sC
;
-------------------------7--w w)R------------------------------------
-
Bumvmhh awR7wR) 
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SR)RR a1 RQ:Rh0R#8F_Do;HO
RSRR RB:hRQR8#0_oDFHSO;
RSRRpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7)ww RR:BbFlFMMC0#RHRk0sC
;
----------------------------7uww-------------------------------------
--
vBmu mhh7aRwRwu
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=4R''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRuRR)  1aQ:Rh0R#8F_Do;HOSR
SRBRRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wuRR:BbFlFMMC0#RHRk0sC
;
-------------------------w-7wRu ---------------------------------------------m
Bvhum Rha7uww RR
RtRR )h Q5BRRR
RRRRRRhRQQ:aRR0LHRR:='R4'
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFHSO;
RSRRRR7:hRQR8#0_oDFH
O;SRRRR u)1R a:hRQR8#0_oDFH
O;SRRRR:B RRQh#_08DHFoO
;SSRRRRiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw wuRB:RFFlbM0CMRRH#0Csk;-

----------------------------7BwwR--------------------------------B

mmvuha hRw7wBR
RR RthQ )B
R5RRRRRRRRQahQRL:RH:0R=jR''R
RR;R2
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFH
O;SRRRR:7RRRQh#_08DHFoOS;
RRRRBqp )RR:Q#hR0D8_FOoH;R
SRBRRp:iRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7BwwRB:RFFlbM0CMRRH#0Csk;R
RR-R
----------------------------7Bww -R------------------------------------------m
Bvhum Rha7Bww RR
RtRR )h Q5BRRR
RRRRRRhRQQ:aRR0LHRR:='Rj'
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFH
O;SRRRR:7RRRQh#_08DHFoOS;
RRRRBqp )RR:Q#hR0D8_FOoH;R
SRBRR Q:Rh0R#8F_Do;HOSR
SRBRRp:iRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Bww RR:BbFlFMMC0#RHRk0sC
;
-------------------------w-7w-hR-----------------------------m
Bvhum Rha7hwwRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=RjR'
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;SS
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:hRRlBFbCFMMH0R#sR0k
C;
----------------7--w whR--------------------------------B-
mmvuha hRw7wh
 RRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''j
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFHSO;
RSRRRR7:hRQR8#0_oDFH
O;SRRRRRB :hRQR8#0_oDFHSO;
RSRRpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww RR:BbFlFMMC0#RHRk0sC
;
-------------------------w7wh-1R--------------------------------
vBmu mhh7aRw1whRR
RR RthQ )BRR5
RRRRRRRRQQhaL:RH:0R=4R''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SR1RR :aRRRQh#_08DHFoO
;SSRRRRiBpRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRw1whRB:RFFlbM0CMRRH#0Csk;-

-------------------------7--w1wh ------------------------------------
--Bumvmhh awR7w h1RR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=R4R'
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SR1RR :aRRRQh#_08DHFoOS;
RRRRBR :Q#hR0D8_FOoH;SS
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w h1RB:RFFlbM0CMRRH#0Csk;-

----------------------------7hww)--------------------------------
--Bumvmhh awR7wRh)
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''R
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HO
RSRR R)1R a:hRQR8#0_oDFHSO;
RSRRpRBiRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww)RR:BbFlFMMC0#RHRk0sCR;
R
RR-------------------------7--w)wh -R----------------------------------
--Bumvmhh awR7w h)RR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=RjR'
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;R
SR7RRRQ:Rh0R#8F_Do;HO
RSRR R)1R a:hRQR8#0_oDFH
O;SRRRR:B RRQh#_08DHFoOS;
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w h)RB:RFFlbM0CMRRH#0Csk;-

-------------------------7--wuwh-------------------------------------
--Bumvmhh awR7wRhu
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=4R''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRuRR)  1aQ:Rh0R#8F_Do;HOSR
SRBRRp:iRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7hwwuRR:BbFlFMMC0#RHRk0sC
;
-------------------------w-7w huR--------------------------------------------B-
mmvuha hRw7whRu 
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=4R''R
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HO
RSRRRR7:hRQR8#0_oDFH
O;SRRRR u)1R a:hRQR8#0_oDFH
O;SRRRR:B RRQh#_08DHFoOS;
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w huRB:RFFlbM0CMRRH#0Csk;-

----------------------------7hwwB-R------------------------------------------B-
mmvuha hRw7wh
BRRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''j
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFH
O;SRRRR:7RRRQh#_08DHFoOS;
RRRRBqp )RR:Q#hR0D8_FOoH;R
SRBRRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:BRRlBFbCFMMH0R#sR0k
C;
----------------------------w-7w hBR-------------------------------------------
vBmu mhh7aRwBwh RR
RtRR )h Q5BRRR
RRRRRRhRQQ:aRR0LHRR:='
j'RRRR2
;SRRRRuam)RS5
RRRRTRR:mRza#_08DHFoO
;SSRRRR:7RRRQh#_08DHFoOS;
RRRRBqp )RR:Q#hR0D8_FOoH;R
SRBRR Q:Rh0R#8F_Do;HOSR
SRBRRp:iRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whRB :FRBlMbFCRM0H0#Rs;kC
-
------------------------------p-7R----------------------------------------
--Bumvmhh apR7RR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=Rj
'RRRRR2
;SRRRRuam)RS5
RRRRTRR:mRza#_08DHFoO
;SSRRRR:7RRRQh#_08DHFoO
;SSRRRR:tRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRR7p:FRBlMbFCRM0H0#Rs;kC
-
----------------------7--p- ----------------------------------m
Bvhum Rha7
p RRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''jRR
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HO
RSRR RB:hRQR8#0_oDFHSO;
RSRRRRt:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7 RR:BbFlFMMC0#RHRk0sC
;
-----------------------------B7pR------------------------------------m
Bvhum Rha7RpB
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRBRRp) qRQ:Rh0R#8F_Do;HOSR
SRtRRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:BRRlBFbCFMMH0R#sR0k
C;
----------------------------p-7B- R---------------------------------
--Bumvmhh apR7B
 RRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''jRR
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HO
RSRRpRB Rq):hRQR8#0_oDFHSO;
RSRRRRt:hRQR8#0_oDFH
O;SRRRR:B RRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRB7p RR:BbFlFMMC0#RHRk0sC
;
-----------------------------u7pR------------------------------------m
Bvhum Rha7Rpu
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=4R''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:#_08DHFoOS;
RRRRu1)  :aRRRQh#_08DHFoO
;SSRRRRRt:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rpu:FRBlMbFCRM0H0#Rs;kC
-
--------------------------7--pRu ------------------------------------
vBmu mhh7aRpRu 
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=4R''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRuRR)  1aRR:Q#hR0D8_FOoH;SS
RRRRtRR:Q#hR0D8_FOoH;R
SRBRR Q:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRu :FRBlMbFCRM0H0#Rs;kC
-
----------------------p-7h-R-----------------------------------------
vBmu mhh7aRp
hRRRRRt  h)RQB5RR
RRRRRQRRhRQa:HRL0=R:R''jRR
RR;R2SR
RRmRu)5aR
RSRRRRT:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HOSR
SRtRRRQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:hRRlBFbCFMMH0R#sR0k
C;
----------------------------p-7h- ----------------------------------m
Bvhum Rha7 phRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=Rj
'RRRRR2
;SRRRRuam)RS5
RRRRTRR:mRza#_08DHFoO
;SSRRRR:7RRRQh#_08DHFoOS;
RRRRBR :Q#hR0D8_FOoH;SS
RRRRtRR:Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7 phRB:RFFlbM0CMRRH#0Csk;R
RR-R
----------------------------7BphR------------------------------------m
Bvhum Rha7BphRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=RjR'
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;R
SR7RRRQ:Rh0R#8F_Do;HO
RSRRpRB Rq):hRQR8#0_oDFH
O;SRRRR:tRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRh7pBRR:BbFlFMMC0#RHRk0sC
;
-----------------------------h7pB- R---------------------------------
--Bumvmhh apR7hRB 
RRRRht  B)QR
5RRRRRRRRRQahQRL:RH:0R=jR''RR
R2RR;RS
RuRRmR)a5R
SRTRRRm:Rz#aR0D8_FOoH;R
SR7RRRQ:Rh0R#8F_Do;HO
RSRRpRB Rq):hRQR8#0_oDFH
O;SRRRR:tRRRQh#_08DHFoOS;
RRRRBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7Bph RR:BbFlFMMC0#RHRk0sC
;
-----------------------------h7pu-R----------------------------------B-
mmvuha hRh7puRR
RtRR )h Q5BRRR
RRRRRRhRQQ:aRR0LHRR:='R4'
RRRRS2;
RRRR)uma
R5SRRRR:TRRamzR8#0_oDFHSO;
RSRRRR7:0R#8F_Do;HO
RSRR)Ru a1 RQ:Rh0R#8F_Do;HOSR
SRtRR:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7h:uRRlBFbCFMMH0R#sR0k
C;
----------------------------p-7hRu ------------------------------------
vBmu mhh7aRp huRR
RR RthQ )BRR5
RRRRRRRRQQhaRR:LRH0:'=R4
'RRRRR2
;SRRRRuam)RS5
RRRRTRR:mRza#_08DHFoO
;SSRRRR:7RRRQh#_08DHFoOS;
RRRRu1)  :aRRRQh#_08DHFoO
;SSRRRR:tRRRQh#_08DHFoOS;
RRRRBR :Q#hR0D8_FOoH
RRRRS2;
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7uph RR:BbFlFMMC0#RHRk0sC
;
--------------------------------)4qvn-14-------------------------m
Bvhum Rha)4qvnR14
RRRRht  B)QR
5RRRRRRRRRQahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jjRj"
RRRR
2;RRRRuam)RS5
SR7m:kRF00R#8F_Do;HO
BSSp:iRRRHM#_08DHFoOS;
S W)RH:RM0R#8F_Do;HO
qSS7RR:H#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
7SSQRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRqnv41:4RRlBFbCFMMH0R#sR0k
C;
--------------------------------v)q4.n1-------------------------B-
mmvuha hRv)q4.n1RR
RR RthQ )BRR5
RRRRRRRRQQhaR_j:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
RRRRRRhRQQ4a_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"RR
R2RR;R
RRmRu)5aR
7SSmRR:FRk0#_08DHFoOC_POs0F584RF0IMF2Rj;S
SBRpi:MRHR8#0_oDFH
O;S)SW RR:H#MR0D8_FOoH;S
Sq:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S7:QRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRqnv41:.RRlBFbCFMMH0R#sR0k
C;RRRR
--------------------------------v)q4cn1-------------------------B-
mmvuha hRv)q4cn1RR
RR RthQ )B
5RRRRRRRRRQahQ_:jRR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RRRRRRRRQQhaR_4:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
RRRRRRhRQQ.a_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R;
RRRRRQRRh_QadRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjjR"
R2RR;R
RRmRu)5aR
7SSmRR:FRk0#_08DHFoOC_POs0F58dRF0IMF2Rj;SR
SiBpRH:RM0R#8F_Do;HO
WSS): RRRHM#_08DHFoOS;
SRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SR7Q:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnR1c:FRBlMbFCRM0H0#Rs;kC
RRRR-
------------------------------q-)v14n7-u4-------------------------m
Bvhum Rha)4qvnu174RR
RtRR )h QRB5
RRRRRRRRQQhaR_j:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jjRR
RR;R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH;S
SBRpi:MRHR8#0_oDFH
O;S)SW RR:H#MR0D8_FOoH;S
SWRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
S7)qRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;SQS7RH:RM0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVqR)v14n7Ru4:FRBlMbFCRM0H0#Rs;kC
-
------------------------------q-)v14n7-u.-------------------------m
Bvhum Rha)4qvnu17.RR
RtRR )h Q5BRRR
RRRRRRhRQQja_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R;
RRRRRQRRh_Qa4RR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjjR"
R2RR;R
RRmRu)5aR
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fs4FR8IFM0R;j2
RSRRpRBiRR:H#MR0D8_FOoH;R
SRWRR): RRRHM#_08DHFoOS;
RRRRWRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
RRRR)Rq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
RRRR7:QRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRqnv41.7uRB:RFFlbM0CMRRH#0Csk;-

-----------------------------)--qnv41c7u-------------------------B-
mmvuha hRv)q47n1u
cRRRRRt  h)RQB5RR
RRRRRQRRh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
";RRRRRRRRQahQ_:4RR0LH_OPC05Fs486RF0IMF2RjRR:=Xj"jj;j"
RRRRRRRRQQhaR_.:HRL0C_POs0F5R468MFI0jFR2=R:RjX"j"jj;R
RRRRRRhRQQda_RL:RHP0_CFO0s654RI8FMR0Fj:2R="RXjjjj"R
RR;R2
RRRR)uma
R5SmS7RF:Rk#0R0D8_FOoH_OPC05FsdFR8IFM0R;j2
BSSp:iRRRHM#_08DHFoOS;
S W)RH:RM0R#8F_Do;HO
WSSq:7RRRHM#_08DHFoOC_POs0F58dRF0IMF2Rj;S
S)Rq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2S;
SR7Q:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4qvnu17cRR:BbFlFMMC0#RHRk0sC
;
--------------------------------)4mvn----------------------------B-
mmvuha hRv)m4
nRRRRRt  h)RQB5RR
RRRRRQRRh_QajRR:L_H0P0COF4s56FR8IFM0RRj2:X=R"jjjj
"RRRRR2R;
RuRRmR)a5S
RRRRR7:mRR0FkR8#0_oDFH
O;SRRRRRq7:MRHR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV)4mvnRR:BbFlFMMC0#RHRk0sC
;
-----------------eQh---------------------------------m
Bvhum RhaQRhe
RRRR)uma
R5RRRRS:mRRamzR8#0_oDFH
O;RRRRS:QRRRQh#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQRhe:FRBlMbFCRM0H0#Rs;kC
-
------------------A--z-wt-------------------------B-
mmvuha hRwAztRR
RuRRm5)a
RRRRRSm:kRF00R#8F_Do;HO
RRRRRSQ:MRHR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRwAztRR:BbFlFMMC0#RHRk0sC
;
-----------------wAz1--------------------m
Bvhum RhaA1zwRR
RRmRu)5aR
RRRRRRRR:mRR0FkR8#0_oDFH
O;RRRRRRRRQRR:H#MR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFAVRzRw1:FRBlMbFCRM0H0#Rs;kC
-
---------------------t-h7----------------
vBmu mhhtaRh
7RRRRRuam)RR5
RSRRtRR:FRk0#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVtRh7:FRBlMbFCRM0H0#Rs;kC
-
------------------e--B-B----------------------B-
mmvuha hRBeBRR
RRmRu)5aR
RRRRRSe:kRF00R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVBReBRR:BbFlFMMC0#RHRk0sC
;
---------------------A-Qz-w----------------------------------
--Bumvmhh aARQz
wRRRRRuam)RR5
RSRRmRR:mRza#_08DHFoOR;
RSRRQRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRARzw:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------mwAz-------------------------------------
--Bumvmhh aARmz
wRRRRRuam)RR5
RSRRmRR:mRza#_08DHFoOR;
RSRRQRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVRARzw:FRBlMbFCRM0H0#Rs;kC
-
----------------------------------A-az-w--------------------------m
Bvhum RhaawAzRR
RRmRu)5aR
RRRRRSm:zRma0R#8F_Do;HO
RRRRRSQ:hRQR8#0_oDFH
O;RRRRShm RQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVARaz:wRRlBFbCFMMH0R#sR0k
C;RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFaVRARzw:FRBlMbFCRM0H"#Rm
";
----------------------------AQmz-w------------------------------B-
mmvuha hRAQmzRw
RuRRmR)a5R
RRmRSRRR:mRzaR0R#8F_Do;HO
RRRRmSQRQ:RhamzR8#0_oDFH
O;RRRRRRSQRQ:RhRRRR8#0_oDFH
O;SRRRRhm RQ:RhRRRR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRAQmz:wRRlBFbCFMMH0R#sR0k
C;
----------------p-ae_71QwAz---------------------------------m
Bvhum Rhaa7pe1A_QzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH;R
RRRRRRARQRQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFReap7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1A_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------eap7m1_A-zw--------------------------------
vBmu mhhaaRp1e7_zmAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRmRRARR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFReap7m1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1A_mz:wRRlBFbCFMMH0R#mR",ARm"
;
-----------------eap7a1_A-zw--------------------------------
vBmu mhhaaRp1e7_zaAwR
RRmRu)5aR
RRRRRSmRm:RzRaR#_08DHFoOR;
RSRRm:ARRamzR0R#8F_Do;HO
RRRRQRSRRR:QRhRR8#0_oDFH
O;SRRRRhm RQ:Rh#RR0D8_FOoH
RRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpRae_71awAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFReap7a1_ARzw:FRBlMbFCRM0H"#Rmm,RA
";
----------------p-ae_71QzmAw--------------------------------B-
mmvuha hReap7Q1_mwAz
RRRR)uma
R5RRRRSRmR:zRma#RR0D8_FOoH;R
RRQRSm:ARRmQhz#aR0D8_FOoH;R
RRRRRRmRQRQ:RhamzR8#0_oDFH
O;RRRRRRSQRQ:Rh0R#8F_Do;HO
RSRR RmhRR:Q#hR0D8_FOoH
RRRR
2;CRM8Bumvmhh aR;
RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpRae_71QzmAwRR:BbFlFMMC0#RHRk0sCR;
RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpRae_71QzmAwRR:BbFlFMMC0#RHRm"Q,mRQA
";
----------------p- e_71QwAz---------------------------------m
Bvhum Rha 7pe1A_QzRw
RuRRm5)a
RRRRRRRR:mRRamzR8#0_oDFH
O;RRRRRRRRQRR:Q#hR0D8_FOoH;R
RRRRRRARQRQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_Qz:wRRlBFbCFMMH0R#QR",ARQ"
;
-----------------e p7m1_A-zw--------------------------------
vBmu mhh aRp1e7_zmAwR
RRmRu)
a5RRRRRRRRmRR:mRza#_08DHFoOR;
RRRRRmRRARR:mRza#_08DHFoOR;
RRRRRQRRRQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7m1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_mz:wRRlBFbCFMMH0R#mR",ARm"
;
-----------------e p7a1_A-zw--------------------------------
vBmu mhh aRp1e7_zaAwR
RRmRu)5aR
RRRRRSmRm:Rz#aR0D8_FOoH;R
RRmRSARR:mRza#_08DHFoOR;
RRRRSRQR:hRQR8#0_oDFH
O;SRRRRhm RQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7a1_ARzw:FRBlMbFCRM0H0#Rs;kC
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_az:wRRlBFbCFMMH0R#mR",ARm"
;
-----------------e p7Q1_mwAz---------------------------------m
Bvhum Rha 7pe1m_QA
zwRRRRuam)RR5
RSRRRRmR:zRma0R#8F_Do;HO
RRRRQSRm:ARRmQhz#aR0D8_FOoH;R
RRRRRRQRRmRR:Qzhma0R#8F_Do;HO
RRRRRRSQ:RRRRQh#_08DHFoOS;
RRRRRhm RQ:Rh0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7Q1_mwAzRB:RFFlbM0CMRRH#0Csk;R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRe p7Q1_mwAzRB:RFFlbM0CMRRH#",QmRAQm"
;

v--Q/uQQRdBHkFLVCRMC08RFCRLRMOFVlHsC
83
--------------------------------7-Q7-)-------------------------
vBmu mhhQaR7R7)
RRRRht  B)QRS5
RRRRTQj_hRQa:HRL0=R:R''j;R
SRTRR4h_QQ:aRR0LHRR:='
j'RRRR2
;SRRRRuam)RS5
RRRRT:jRRamzR8#0_oDFH
O;SRRRRRT4:zRma0R#8F_Do;HOSR
SR7RRRQ:Rh0R#8F_Do;HO
RSRRpRBiQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7R7):FRBlMbFCRM0H0#Rs;kC
-
------------------------------Q--7B7)-------------------------
--Bumvmhh a7RQ7R)B
RRRRht  B)QR
5RSRRRR_TjQahQRL:RH:0R=jR''S;
RRRRTQ4_hRQa:HRL0=R:R''j
RRRRS2;
RRRR)uma
R5SRRRRRTj:zRma0R#8F_Do;HO
RSRR4RTRm:Rz#aR0D8_FOoH;SS
RRRR7RR:Q#hR0D8_FOoH;R
SRBRRp) q:hRQR8#0_oDFHSO;
RSRRpRBiQ:Rh0R#8F_Do
HORRRR2
;SCRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7B7)RB:RFFlbM0CMRRH#0Csk;-

-------------------------Q--7_7)v- v---------------------------------
--Bumvmhh a7RQ7v)_ 
vRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"S
2;S)uma
R5SjSTRF:Rk#0R0D8_FOoH;SS
SRT4:kRF00R#8F_Do;HOSS
S7RR:H#MR0D8_FOoH;S
SQiBpRH:RM0R#8F_Do;HO
uSSBRpi:MRHR8#0_oDFH
O;S S)1R a:MRHR8#0_oDFH
O;SqSW7R7):MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RSRR)7q7)RR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R
j2S
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7_7)vR v:FRBlMbFCRM0H0#Rs;kC
-
------------------------------7m7)--------------------
--Bumvmhh a7Rm7
)RRRRRt  h)RQB5RR
RRRRRaRRXiBp_pumRL:RH:0R=jR''-;R-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bkRRRRRRRR
RRRRRRRRhBm1haqahRQQ:aRR8#0_oDFH:OR=jR''RR
R2RR;RS
RuRRmR)a5SR
RRRRT:jRRamzR8#0_oDFHSO;
RSRR4RTRm:Rz#aR0D8_FOoH;SS
RRRR7:jRRRQh#_08DHFoOS;
RRRR7:4RRRQh#_08DHFoOS;
RRRRa:XRRRQh#_08DHFoOS;
RRRRBRpi:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7Rm7:)RRlBFbCFMMH0R#sR0k
C;
-------------------------------m)77B--------------------
--Bumvmhh a7Rm7R)B
RRRRht  B)QR
5RRRRRRRRRapXBim_upRR:LRH0:'=RjR';-j-''H:)#oHMRoC8CkRF00bk;4R''N:wDMDHo8RCoFCRkk0b0R
RRRRRRmRBhq1ahQaRhRQa:0R#8F_DoRHO:'=RjR'
R2RR;R
RRmRu)5aR
RSRRjRTRm:Rz#aR0D8_FOoH;R
SRTRR4RR:mRza#_08DHFoOS;
RRRR7:jRRRQh#_08DHFoOS;
RRRR7:4RRRQh#_08DHFoOS;
RRRRa:XRRRQh#_08DHFoOS;
RRRRBRpi:hRQR8#0_oDFH
O;SRRRR Bpq:)RRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7m7):BRRlBFbCFMMH0R#sR0k
C;
----------------------------7m7) _vv------------------------------------m
Bvhum Rham)77_vv RR
RR RthQ )BS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k;C"
RRRRRRRRBaXpui_m:pRR0LHRR:=';j'R'--j)':HM#Ho8RCoFCRkk0b0';R4w':NHDDMCoR8RoCFbk0kR0
RRRRRaRRB_pi1)mzB: RRs#0HRMo:"=R7WT1"R
RR;R2
RRRR)uma
R5STSRjRR:FRk0#_08DHFoO
;SSTSR4RR:FRk0#_08DHFoO
;SSaSRBRpi:MRHR8#0_oDFH
O;SuSRBRpi:MRHR8#0_oDFH
O;S)SR a1 RH:RM0R#8F_Do;HO
RSS7:jRRRHM#_08DHFoOS;
S4R7RH:RM0R#8F_Do;HO
RSSa:XRRRHM#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)77_vv RB:RFFlbM0CMRRH#0Csk;-

----------------------------------------Q17 c-------------------------------
vBmu mhhQaR7c 1Rt
S )h Q5BR
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)h:RRRs#0HRMo:"=R0Csk"2
S;u
SmR)a5S
S7RR:Q#hR0D8_FOoH;S
SBQqpARR:Q#hR0D8_FOoH;S
S)  1aRR:Q#hR0D8_FOoH;S
SwiBpRQ:Rh0R#8F_Do;HO
uSSBRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ R1c:FRBlMbFCRM0H0#Rs;kC
-
-------------------------Q17 c _vv--------------------------------
--Bumvmhh a7RQ _1cvR v
CSoMHCsOS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"S
2;S)umaS5
S)7, a1 RQ:Rh0R#8F_Do;HO
BSSqApQRQ:Rh0R#8F_Do;HO
QSSB,piwiBp,puBiRR:Q#hR0D8_FOoH;S
SW7q7)RR:Q#hR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
)SSq)77RQ:Rh0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFHSO
R
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVR7c 1_vv RB:RFFlbM0CMRRH#0Csk;-

---------------------------------Q--e Q7m-------------------------------
vBmu mhhQaRe Q7mRR
RtRR )h Q5BR
tSS1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)h:RRRs#0HRMo:"=R0Csk"R
RR;R2
RRRR)uma
R5SRS7:hRQR8#0_oDFH
O;S S)1R a:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;SBSwp:iRRRQh#_08DHFoOS;
SpuBiRR:Q#hR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH;S
ST:.RRamzR8#0_oDFH
O;SdSTRm:Rz#aR0D8_FOoH;S
ST:cRRamzR8#0_oDFH
O;S6STRm:Rz#aR0D8_FOoH;S
ST:nRRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRQQe7R m:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------- Q71-U----------------------------------
--Bumvmhh a7RQ R1U
RRRRht  B)QRS5
RRRRt 1)hRR:#H0sM:oR=VR"NCD#"S;
S)p1 RhR:0R#soHMRR:="k0sCR"
R2RR;R
RRmRu)5aR
7SS,1)  :aRRRQh#_08DHFoOS;
SpBqQ:ARRRQh#_08DHFoOS;
SpwBiB,up:iRRRQh#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoOS;
SRT.:zRma0R#8F_Do;HO
TSSdRR:mRza#_08DHFoOS;
SRTc:zRma0R#8F_Do;HO
TSS6RR:mRza#_08DHFoOS;
SRTn:zRma0R#8F_Do;HO
TSS(RR:mRza#_08DHFoOR
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 URR:BbFlFMMC0#RHRk0sC
;
------------------------- Q71vU_ -v--------------------------B-
mmvuha hR Q71vU_ 
vRRRRRt  h)RQB5R
SRtRR1h) R#:R0MsHo=R:RN"VD"#C;S
Sp 1)h:RRRs#0HRMo:"=R0Csk"R
RR;R2
RRRR)uma
R5S,S7)  1aRR:Q#hR0D8_FOoH;S
SBQqpARR:Q#hR0D8_FOoH;S
SwiBp,pQBiB,up:iRRRQh#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoOS;
SRT.:zRma0R#8F_Do;HO
TSSdRR:mRza#_08DHFoOS;
SRTc:zRma0R#8F_Do;HO
TSS6RR:mRza#_08DHFoOS;
SRTn:zRma0R#8F_Do;HO
TSS(RR:mRza#_08DHFoOS;
S7Wq7:)RRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;S
S)7q7)RR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ _1UvR v:FRBlMbFCRM0H0#Rs;kC
-
-------------------------------------Q17 4-j---------------------------------
vBmu mhhQaR74 1jRR
RtRR )h Q5BR
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
pSS1h) RRR:#H0sM:oR=0R"s"kC
RRRR
2;RRRRuam)RS5
S)7, a1 RQ:Rh0R#8F_Do;HO
BSSqApQRQ:Rh0R#8F_Do;HO
wSSB,piuiBpRQ:Rh0R#8F_Do;HO
TSSjRR:mRza#_08DHFoOS;
SRT4:zRma0R#8F_Do;HO
TSS.RR:mRza#_08DHFoOS;
SRTd:zRma0R#8F_Do;HO
TSScRR:mRza#_08DHFoOS;
SRT6:zRma0R#8F_Do;HO
TSSnRR:mRza#_08DHFoOS;
SRT(:zRma0R#8F_Do;HO
TSSURR:mRza#_08DHFoOS;
SRTg:zRma0R#8F_Do
HORRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ j14RB:RFFlbM0CMRRH#0Csk;-

---------------------------------7-Q n14-------------------------------------m
Bvhum RhaQ17 4Rn
RtRR )h Q5BR
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k
C"RRRR2R;
RuRRmR)a5S
S7 ,)1R a:hRQR8#0_oDFH
O;SqSBpRQA:hRQR8#0_oDFH
O;SBSwpui,BRpi:hRQR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFH
O;S.STRm:Rz#aR0D8_FOoH;S
ST:dRRamzR8#0_oDFH
O;ScSTRm:Rz#aR0D8_FOoH;S
ST:6RRamzR8#0_oDFH
O;SnSTRm:Rz#aR0D8_FOoH;S
ST:(RRamzR8#0_oDFH
O;RRRRRRRRT:URRamzR8#0_oDFH
O;SgSTRm:Rz#aR0D8_FOoH;S
STR4j:zRma0R#8F_Do;HO
TSS4:4RRamzR8#0_oDFH
O;S4ST.RR:mRza#_08DHFoOS;
SdT4Rm:Rz#aR0D8_FOoH;S
STR4c:zRma0R#8F_Do;HO
TSS4:6RRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71R4n:FRBlMbFCRM0H0#Rs;kC
-
----------------------m--1c )-----------------------------B-
mmvuha hR m1)
cRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sC
";RRRRRRRR]RWp:0R#soHMRR:="DVN#;C"R"--0Csk"";RV#NDCR"
RRRRRaRRXiBp_pumRL:RH:0R=jR''-R-':j')HH#MCoR8RoCFbk0kR0;':4'wDNDHRMoCC8oR0Fkb
k0S
2;S)uma
R5SjS7RH:RM0R#8F_Do;HO
7SS4RR:H#MR0D8_FOoH;S
S7:.RRRHM#_08DHFoOS;
SR7d:MRHR8#0_oDFH
O;SXSajRR:H#MR0D8_FOoH;S
SaRX4:MRHR8#0_oDFH
O;SBSup:iRRRHM#_08DHFoOS;
S1)  :aRRRHM#_08DHFoOS;
SpwBiRR:H#MR0D8_FOoH;S
ST:jRRamzR8#0_oDFH
O;S4STRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 cRR:BbFlFMMC0#RHRk0sC
;
----------------- m1)vc_ -v------------------------------B-
mmvuha hR m1)vc_ 
vRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sC
";SWS]pRR:#H0sM:oR=VR"NCD#"R;
RRRRRaRRXiBp_pumRL:RH:0R=jR''-;-':j')HH#MCoR8RoCFbk0kR0;':4'wDNDHRMoCC8oR0Fkb
k0RRRRRRRRaiBp_z1m)RB :0R#soHMRR:="17TWR"RRSR
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SjaXRH:RM0R#8F_Do;HO
aSSX:4RRRHM#_08DHFoOS;
SpuBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SwiBpRH:RM0R#8F_Do;HO
aSSBRpi:MRHR8#0_oDFH
O;SjSTRm:Rz#aR0D8_FOoH;S
ST:4RRamzR8#0_oDFHSO
2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rm _)cvR v:FRBlMbFCRM0H0#Rs;kC
-
------------------e-mQm7 ---------------------------------B-
mmvuha hRQme7R m
 SthQ )BS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sCS"
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SR7c:MRHR8#0_oDFH
O;S6S7RH:RM0R#8F_Do;HO
7SSnRR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SRST:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVRe Q7mRR:BbFlFMMC0#RHRk0sC
;
--------------------m)1 U-----------------------------------
vBmu mhhmaR1U )RR
RR RthQ )B
R5RRRRS)t1 :hRRs#0HRMo:"=RV#NDC
";RRRRS)p1 :hRRs#0HRMo:"=R0Csk"R;
RRRRR]RRW:pRRs#0HRMo:"=RV#NDC
";RRRRRRRRapXBim_upRR:LRH0:'=Rj-'R-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bk
RRRR
2;RRRRuam)RR5
RRRRR7RSjRR:H#MR0D8_FOoH;R
RRRRRR4S7RH:RM0R#8F_Do;HO
RRRRRRRSR7.:MRHR8#0_oDFH
O;RRRRRSRR7:dRRRHM#_08DHFoOR;
RRRRR7RScRR:H#MR0D8_FOoH;R
RRRRRSR76:MRHR8#0_oDFH
O;RRRRRSRR7:nRRRHM#_08DHFoOR;
RRRRR7RS(RR:H#MR0D8_FOoH;R
RRRRRRXSajRR:H#MR0D8_FOoH;R
RRaRSX:4RRRHM#_08DHFoOS;
RRRRaRX.:MRHR8#0_oDFH
O;SRRRRdaXRH:RM0R#8F_Do;HO
RSRRBRup:iRRRHM#_08DHFoOS;
RRRR)  1aRR:H#MR0D8_FOoH;R
SRwRRBRpi:MRHR8#0_oDFH
O;RRRRRSRRT:jRRamzR8#0_oDFH
O;RRRRRSRRT:4RRamzR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1):URRlBFbCFMMH0R#sR0k
C;
----------------1-m _)Uv- v-----------------------------
--Bumvmhh a1Rm _)UvR v
 SthQ )BS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sC
";SWS]pRR:#H0sM:oR=VR"NCD#"R;
RRRRRaRRXiBp_pumRL:RH:0R=jR''R;
RRRRRaRRB_pi1)mzB: RRs#0HRMo:"=R7WT1"2
S;u
SmR)a5S
S7:jRRRHM#_08DHFoOS;
SR74:MRHR8#0_oDFH
O;S.S7RH:RM0R#8F_Do;HO
7SSdRR:H#MR0D8_FOoH;S
S7:cRRRHM#_08DHFoOS;
SR76:MRHR8#0_oDFH
O;SnS7RH:RM0R#8F_Do;HO
7SS(RR:H#MR0D8_FOoH;S
SaRXj:MRHR8#0_oDFH
O;SXSa4RR:H#MR0D8_FOoH;S
SaRX.:MRHR8#0_oDFH
O;SXSadRR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SBSap:iRRRHM#_08DHFoOS;
SRTj:zRma0R#8F_Do;HO
TSS4RR:mRza#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR m1)vU_ :vRRlBFbCFMMH0R#sR0k
C;
-------------------- m1)-4j---------------------------------B-
mmvuha hR m1)R4j
 SthQ )B
R5S1St)R h:0R#soHMRR:="DVN#;C"
pSS1h) R#:R0MsHo=R:Rs"0k
C"S
2;S)uma
R5SjS7RH:RM0R#8F_Do;HO
7SS4RR:H#MR0D8_FOoH;S
S7:.RRRHM#_08DHFoOS;
SR7d:MRHR8#0_oDFH
O;ScS7RH:RM0R#8F_Do;HO
7SS6RR:H#MR0D8_FOoH;S
S7:nRRRHM#_08DHFoOS;
SR7(:MRHR8#0_oDFH
O;SUS7RH:RM0R#8F_Do;HO
7SSgRR:H#MR0D8_FOoH;S
SuiBpRH:RM0R#8F_Do;HO
)SS a1 RH:RM0R#8F_Do;HO
wSSBRpi:MRHR8#0_oDFH
O;SRST:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR14 )jRR:BbFlFMMC0#RHRk0sC
;
--------------------m)1 4-n----------------------------------m
Bvhum Rham)1 4
nRSht  B)QRS5
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R h:0R#soHMRR:="k0sCS"
2S;
uam)RS5
SR7j:MRHR8#0_oDFH
O;S4S7RH:RM0R#8F_Do;HO
7SS.RR:H#MR0D8_FOoH;S
S7:dRRRHM#_08DHFoOS;
SR7c:MRHR8#0_oDFH
O;S6S7RH:RM0R#8F_Do;HO
7SSnRR:H#MR0D8_FOoH;S
S7:(RRRHM#_08DHFoOS;
SR7U:MRHR8#0_oDFH
O;SgS7RH:RM0R#8F_Do;HO
RRRRRRRRj74RH:RM0R#8F_Do;HO
7SS4:4RRRHM#_08DHFoOS;
S.74RH:RM0R#8F_Do;HO
7SS4:dRRRHM#_08DHFoOS;
Sc74RH:RM0R#8F_Do;HO
7SS4:6RRRHM#_08DHFoOS;
SpuBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SwiBpRH:RM0R#8F_Do;HO
TSSRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVm)1 4:nRRlBFbCFMMH0R#sR0k
C;
--------------------7Qm Ypq---------------------------------
--
vBmu mhhQaRmp7 q
YRSht  B)QRR5R
RRRRRRRR1B_aQqaBp_7YRR:HCM0oRCs:j=RRR--j.~4(R
RR;R2RR
RRmRu)5aR
7SSQRR:Q#hR0D8_FOoH;S
S1q7auRR:Q#hR0D8_FOoH;S
S1h aRQ:Rh0R#8F_Do;HO
eSSq pzRQ:Rh0R#8F_Do;HO
7SSmRR:mRza#_08DHFoOS;
SR7w:zRma0R#8F_Do
HOS
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFQVRmp7 q:YRRlBFbCFMMH0R#sR0k
C;
--------------------vQ ---------------------------------B-
mmvuha hRvQ Rt
S )h Q
B5SQSWhZ1Q RR:#H0sM:oR=1R"vpqp"S;
S)t1 :hRRs#0HRMo:"=RV#NDC
";S1Sp)R hR#:R0MsHo=R:Rs"0k
C"S
2;S)uma
R5SRS7:MRHR8#0_oDFH
O;SpSBiRR:H#MR0D8_FOoH;S
S)  1aRR:H#MR0D8_FOoH;S
SviBp:MRHR8#0_oDFH
O;SqSptRR:FRk0#_08DHFoOS;
Sqp 7RR:FRk0#_08DHFoO2
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRvQ RB:RFFlbM0CMRRH#0Csk;-

-----------------------------B--pQi7e------------------------
--Bumvmhh apRBie7Q
RRRRht  B)Q5R
SRRRR7_Qev m7R1:Rah)Qt=R:R"".;-R-R"".,dR"3,6"R""c,6R""",RUS"
RRRRR)t1 :hRR)1aQRht:"=RV#NDC-"R-VR"NCD#"",R0Csk"R
SR2RR;R
RRmRu)
a5RRRRRRRRRp]BiRQh:hRQR8#0_oDFH
O;SRRRR R)1h aRQ:Rh0R#8F_Do;HO
RSRRBRRqApQRQ:RM0R#8F_Do;HO
RSRRBRRpzimaRR:mRza#_08DHFoOR
RRRRRR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFVB7piQ:eRRlBFbCFMMH0R#sR0k
C;
--------------------------------B7] -h----------------------------------
--Bumvmhh a]R7B
 hRRRRuam)RS5
RiBpmRza:zRma0R#8F_Do;HOSR
SB: RRRQh#_08DHFoO
;SSpRBiRQh:hRQR8#0_oDFHRO
R2RR;CS
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV]R7BR h:FRBlMbFCRM0H0#Rs;kCRRRR
-
--------------7--T-1------------------------------
--Bumvmhh aTR71R
RR RthQ )BS5
RRRRwmQw_7vm  _1pRR:LRH0:'=Rj-';-QRwwlmRFR8C#CCDOR0:',j'7R7)lFClsl$RF;8C':4'R7t7)FRl8SC
S_)7u)haRL:RHP0_CFO0s=R:Rj"jj-";-wwQmCRsNb8RF0HMC#sRCH00MSo
S17T_7vm RR:#H0sM:oR=XR"4R";-"-RX,4""_X.7.7)"X,".7_7),d"""Xc,."X_)77dX_ aR"
RRRRR]RRW:pRRs#0HRMo:"=RV#NDC-";-s"0k;C"RN"VD"#C
RRRR1St)R h:0R#soHMRR:="DVN#RC"-N-VD,#CRk0sC2
S;R
RRmRu)
a5RRRRRRRR7QT1hB,upwi,B,pi)  1aRR:H#MR0D8_FOoH;S
S)7 qRH:RM0R#8F_Do_HOP0COFds5RI8FMR0Fj
2;SBS)p i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
7SSpap1 Wu,1ua RH:RM0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;SpS)mhq7,vR)m,e RQ)7)],RmRp7:MRHR8#0_oDFH
O;RRRRRRRRWqpm7Rh,Wevm W,R7RQ):MRHR8#0_oDFH
O;RRRRRRRR7)T1gRj,7WT1j7,RT.1W(:jRR0FkR8#0_oDFH
O;SuS)maQh,uRWmaQhRF:Rk#0R0D8_FOoH_OPC05Fs.FR8IFM0R;j2
)SSeQqp7A,)za)1,wR)p,qtRpWwq:tRR0FkR8#0_oDFHRO
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR17TRB:RFFlbM0CMRRH#0Csk;-

----------------7-pp--------------------------------
vBmu mhh7aRpRp
RtRR )h Q
B5RRRRRRRR7_ppwBm) RR:HCM0oRCs:j=R;4--:FRVsROCD	FOR8NMR8OFCj;R:FRO8DC/FRO	oCCMsCN08sRVF7lRpDpRF
FbRRRRRRRR7_Qe1R p:HRL0=R:R''4;j--,sMFlRNDD	FOR8lFC4;R,#VN0FRDOl	RF
8CSRRRR7Bm q1BpRR:1Qa)h:tR=jR"j;j"-j-j44Rjj4Rj4jR4jjR444R4j4R44R
RRRRRRBR1q p_hRR:1Qa)h:tR=0R"s"kC-s-0kVC,NCD#
RRRR
2;RRRRuam)5R
RRRRRRpRBi:QhQ#hR0D8_FOoH:j=''R;
RRRRR1RRa:muRRQM#_08DHFoO':=j
';RRRRRRRR)  1aRR:Q#MR0D8_FOoH:j=''R;
RRRRRzRRuB7hhRap:MRQR8#0_oDFH=O:';j'
RRRRRRRRBpmiRR:mRza#_08DHFoOR;
RRRRR1RRaR u:zRma0R#8F_Do_HOP0COF(s5RI8FMR0FjR2
RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7pRR:BbFlFMMC0#RHRk0sC
;
-----------------------------p-7pY7p-------------------------------------
--Bumvmhh apR7pY7p
RRRRht  B)Q5R
RRRRRRpR7ph_Q1R p:HRL0=R:R''j;-R-':j'LN$b#l#RF,8CR''4:#RkCDR8DC_8DRN$ODCD
RRRRRRRRY7p_t1QhRR:LRH0:'=RjR';-'-Rj'':+R',R''4:-R''R
RRRRRRpR7Y7_qKRR:HCM0oRCs:j=RRj--~6.6,DR8$H_#ojM=RD:8$8_N[8;RD#$_H=oM4-:R.+6n8_D$N
8[RRRR2R;
RuRRm5)a
RRRRRRRRp7p1ua RQ:Rh0R#8F_Do_HOP0COF(s5RI8FMR0Fj
2;RRRRRRRRBQpihh:QR8#0_oDFH
O;RRRRRRRR7,Q)p7mqhm,veR :Q#MR0D8_FOoH;R
RRRRRRpRBiamzRm:Rz#aR0D8_FOoH;R
RRRRRRpRwq:tRRamzR8#0_oDFHRO
RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7pY7pRB:RFFlbM0CMRRH#0Csk;-

-----------------Bm1_adq----------------------------
vBmu mhhmaR1dB_q
aRRRRRt  h)RQB5R
RRRRRR)Rw 7T_Q:eRR0HMCsoCRR:=4RjjR.--~U4.,DFM$PRCCMMRkRl
R2RR;R
RRmRu)5aR
RSRR1RmBamzRF:Rk#0R0D8_FOoH
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFmVR1dB_q:aRRlBFbCFMMH0R#sR0k
C;RRRR
--------------------------------17B-------------------------------------m
Bvhum Rha7
B1RRRRt  h)RQB5S
S7_B1v m7R#:R0MsHo=R:RQ")1tQh"RRR-p-BiBj,p,i4B.pi,iBpdh,t7B,eBQ,)1tQh,pwqptQh,iBpjh_t7p,Biej_BBB,p_i4t,h7B4pi_BeB,iBp.h_t7p,Bie._BBB,p_idt,h7Bdpi_BeB
;S2
mSu)5aR
BSSpRij:hRQR8#0_oDFH
O;SpSBi:4RRRQh#_08DHFoOS;
SiBp.RR:Q#hR0D8_FOoH;S
SBdpiRQ:Rh0R#8F_Do;HO
BSSp i1pRR:Q#hR0D8_FOoH_OPC05FsdFR8IFM0R;j2
1SS mpw)RB :hRQR8#0_oDFH
O;SpSBiamzRm:Rz#aR0D8_FOoH
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV7RB1:FRBlMbFCRM0H0#Rs;kCRRRR
-
------------------------------T-7B- ----------------------------------
--Bumvmhh aTR7BR 
RuRRmR)a5R
SBmpiz:aRRamzR8#0_oDFHSO;
BSR RR:Q#hR0D8_FOoH;SS
RiBpQ:hRRRQh#_08DHFoOR
RR;R2SM
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRB7T RR:BbFlFMMC0#RHRk0sCR;RRRR
R-R
---------------------m-)v----------------------------m
Bvhum Rha)Rmv
RRRRht  B)QR
5RSQRAaQ_W7Ra]:MRH0CCos=R:4
;SS R)qv7_mR7 :HRL0=R:R''j;R
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRRRRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiB,R B,m  ,)1, aWR) :MRHR8#0_oDFH
O;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRv)mRB:RFFlbM0CMRRH#0Csk;-
-----------------------------)Xmvg-R------------------------------------------
--Bumvmhh amR)vRXg
RRRRht  B)QR
5RRRRRA_QaWaQ7]RR:HCM0oRCs:;=g
RRRRq) 7m_v7: RR0LHR':=j
';RRRRA_pi1R p:HRL0C_POs0FRR:="jjj"R;
R)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBRRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
R
RRRR2R;
RuRRmR)a5R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
BSRpRi,Bm ,B) , a1 , W)RH:RM0R#8F_Do;HO
RRRRASRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
qSR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF)VRmgvXRB:RFFlbM0CMRRH#0Csk;-

-----------------u-1-------------------------------------
--Bumvmhh auR1RR
RR RthQ )B
R5SQRAaQ_W7Ra]:MRH0CCos=R:dR.;-4-R,,R.RRc,U4,Rnd,R.R
S)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS)RWQ_a v m7RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiB,R B,m  ,)1, aWR) :MRHR8#0_oDFH
O;S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds54FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR1RB:RFFlbM0CMRRH#0Csk;-

-------------------------1--u-Xg-------------------------------------B-
mmvuha hRX1ugRR
RtRR )h Q5BRRR
SA_QaWaQ7]RR:HCM0oRCs:;=g
)SR _q7v m7RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
RQW)av _mR7 :HRL0C_POs0FR":=j;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;R
SB,piR,B m,B )  1a),W RR:H#MR0D8_FOoH;R
Sq:7RRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
RR7Q:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2R

R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRX1ugRR:BbFlFMMC0#RHRk0sC
;




---------------------------------7-1u-A--------------------------------------m
Bvhum Rha1A7uRR
RR RthQ )BRR5
RSRRQRAaQ_W7_a]jRR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.SRRRRaAQ_7WQa4]_RH:RMo0CC:sR=;4nRR--4.,R,,RcRRU,4Rn,dS.
RRRR)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CRRRRRRRRA_pi1_ pjRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRRiAp_p1 _:4RR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SRBRRp,iqBApi, RBq ,BAB,m  ,)1q a,1)  RaA:MRHR8#0_oDFH
O;SRRRRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRRRRRiAp1q p,iAp1A pRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SRRRRR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu17ARR:BbFlFMMC0#RHRk0sC
;
---------------------------------7-1uAXg-------------------------------------
--Bumvmhh a7R1uAXgRR
RR RthQ )BRR5
RSRRQRAaQ_W7_a]jRR:HCM0oRCs:U=4;-R-RRg,4RU,dSn
RRRRA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4,nRd
RSRR R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SRARRp1i_ jp_RL:RHP0_CFO0s=R:Rj"jj
";SRRRRiAp_p1 _:4RR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
RRRRRR2R;
RuRRmR)a5R
SR7RRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;SRRRRiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 ARR:H#MR0D8_FOoH;R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRRARRp i1pAq,p i1p:ARRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SR7RRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF1VR7guXARR:BbFlFMMC0#RHRk0sC
;
----------------------------7-uA-------------------------------------
-
Bumvmhh auR7ARR
RtRR )h Q5BR
RSSA_QaWaQ7]R_j:MRH0CCos=R:4Rn;
RSSA_QaWaQ7]R_4:MRH0CCos=R:4Rn;
RSS)7 q_7vm :jRR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
RSS)7 q_7vm :4RR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
RSSWa)Q m_v7R j:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RSSWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RRRRASRp1i_ jp_RL:RHP0_CFO0s=R:Rj"jj
";RRRRSpRAi _1pR_4:HRL0C_POs0FRR:="jjj"R;
RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSSQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSSQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
j"RRRR2R;
RuRRmR)a5S
SRq7m,A7mRF:Rk#0R0D8_FOoH_OPC05Fs486RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,42S;
SpRBiBq,p,iARqB ,AB , mBqB,m )A, a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
RRRRSA1pi ,pqA1pi RpA:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRu:ARRlBFbCFMMH0R#sR0k
C;
----------------------------X7ug-A--------------------------------------m
Bvhum Rha7guXARR
RtRR )h Q5BRRR
SRARRQWa_Q]7a_:jRR0HMCsoCR4:=U-;R-,RgR
4USRRRRaAQ_7WQa4]_RH:RMo0CC:sR=;4URR--g4,RUR
SR)RR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CSRRRRq) 7m_v7R 4:HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SRWRR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8CSRRRRQW)av _m47 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
RRRRRRpRAi _1pR_j:HRL0C_POs0FRR:="jjj"R;
RRRRRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
RSRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
RRRR
2;RRRRuam)RS5
RRRR7,mq7RmA:kRF00R#8F_Do_HOP0COF4s5(FR8IFM0RRj2:O=RF_MP#_08DHFoOC_POs0F54j,U
2;SRRRRiBpqp,BiRA,B, qB, AmqB , mBA ,)1q a,1)  ,aAWq) , W)ARR:H#MR0D8_FOoH;R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2S;
RRRR7RQq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;RRRRRRRRA1pi ,pqA1pi RpA:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RRRR7RQA:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRX7ug:ARRlBFbCFMMH0R#sR0k
C;




--------------------------------1--7-u--------------------------------------m
Bvhum Rha1R7u
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
S7:QRRRHM#_08DHFoOC_POs0F5Rd48MFI0jFR2R
RR;R2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV1R7u:FRBlMbFCRM0H0#Rs;kC
-
---------------------------------1X7ug---------------------------------------
vBmu mhh1aR7guXRR
RR RthQ )BRR5
ASRQWa_Q]7a_:jRR0HMCsoCR4:=U-;R-,RgR,4UR
dnSQRAaQ_W7_a]4RR:HCM0oRCs:U=4;-R-RRg,4RU,dSn
Rq) 7m_v7: RR0LHRR:=';j'RR--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
ASRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRRR
RRRR
2;RRRRuam)RS5
RR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;R
SBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoOS;
Rqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV7R1uRXg:FRBlMbFCRM0H0#Rs;kC
-S
---------------------------------7s1u---------------------------------------
vBmu mhhsaR1R7u
RRRRht  B)QR
5RSQRAaQ_W7_a]jRR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;-R-RR4,.c,R,,RUR,4nR
d.S R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hBShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRR
R2RR;R
RRmRu)5aR
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1a:ARRRHM#_08DHFoOS;
Rqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;SQR7RH:RM0R#8F_Do_HOP0COFds54FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rs7:uRRlBFbCFMMH0R#sR0k
C;
--------------------------------s--1X7ug---------------------------------------
vBmu mhhsaR1X7ugRR
RtRR )h Q5BRRR
SA_QaWaQ7]R_j:MRH0CCos=R:4RU;-g-R,UR4,nRd
ASRQWa_Q]7a_:4RR0HMCsoCR4:=U-;R-,RgR,4UR
dnS R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCR
SA_pi1R p:HRL0C_POs0FRR:="jjj"R;
RRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;R-h1YBq,R1BYh
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRRR
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 ARR:H#MR0D8_FOoH;R
Sq,7qqR7A:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RR7Q:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFR7s1uRXg:FRBlMbFCRM0H0#Rs;kC




-
----------------------mb)v----------------------------m
Bvhum Rhabv)mRR
RR RthQ )BRR5
RSRRQRAaQ_W7Ra]:MRH0CCos=R:4
;SSRRRRq) 7m_v7: RR0LHRR:=';j'
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
SRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRRRR
RRRR
2;RRRRuam)RS5
RRRR7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
RSRRpRBiB,R m,RBR ,)  1aRR:H#MR0D8_FOoH;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFbVR)Rmv:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------bv)mX-gR--------------------------------------------
vBmu mhhbaR)XmvgRR
RtRR )h Q5BRRR
RRRRRRQRAaQ_W7Ra]:MRH0CCos=R:gR;
RRRRR)RR _q7v m7RL:RH:0R=''j;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hRB
RRRRRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRRR

R2RR;R
RRmRu)5aR
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RRRRB,piR,B R mB, R)1R a:MRHR8#0_oDFH
O;SRRRRRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2
R2RR;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRmb)vRXg:FRBlMbFCRM0H0#Rs;kC



---------------------s--)-mv-------------------------
--Bumvmhh a)Rsm
vRRRRRt  h)RQB5SR
RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SR
SR)RR _q7v m7RL:RH:0R=jR''R;
RRRRRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRRRRR
RR;R2
RRRR)uma
R5SRRRRR7m:kRF00R#8F_Do_HOP0COFds54FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2d.;R
SRBRRpRi,BR ,m,B R1)  :aRRRHM#_08DHFoOR;
RSRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGFsVR)Rmv:FRBlMbFCRM0H0#Rs;kC
-
-----------------------------sv)mX-gR--------------------------------------------
vBmu mhhsaR)XmvgRR
RtRR )h Q5BRRR
RRRRRRQRAaQ_W7Ra]:MRH0CCos=R:gR;
RRRRR)RR _q7v m7RL:RH:0R=''j;R
RRRRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBR
RRRRRRhRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR
R
RR;R2
RRRR)uma
R5SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2S;
RiBp, RB,BRm ),R a1 RH:RM0R#8F_Do;HO
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRV)RsmgvXRB:RFFlbM0CMRRH#0Csk;

S
-----------------------------7u-------------------------------------B-
mmvuha hRR7u
RRRRht  B)QRS5
SQRAaQ_W7_a]jRR:HCM0oRCs:n=4;SR
SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;SR
S R)qv7_mj7 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
S)RWQ_a v m7jRR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8SC
S)RWQ_a v m74RR:L_H0P0COF:sR=jR"jR";-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8RC
RSRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";RRRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBS
SRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S
SRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj
RRRR
2;RRRRuam)RS5
SmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R468MFI0jFR2O:=F_MP#_08DHFoOC_POs0F54j,n
2;SBSRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;SqSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2R;
RSRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
RRRR
2;CRM8Bumvmhh aS;
Ns00H0LkC$R#MD_LN_O	LRFGF7VRuRR:BbFlFMMC0#RHRk0sC
;
----------------------------7guX-------------------------------------
--Bumvmhh auR7X
gRRRRRt  h)RQB5SR
RaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUR
SA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4
)SR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8CS R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8SC
RQW)av _mj7 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCR
SWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
RRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1hSB
RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"S;
RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRR
R2RR;R
RRmRu)5aR
7SRm7q,m:ARR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5j4;U2
BSRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R
S7RQq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2S;
RA7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R
j2RRRR2C;
MB8Rmmvuha h;N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR7X:gRRlBFbCFMMH0R#sR0k
C;
----------------------------u7164n_..X41-zv-------------------------------------B-
mmvuha hRu7164n_..X41
zvRRRRoCCMs5HO
qSSjt) _iBpR#:R0MsHo=R:RY"Au1q1"-;R-AR"Y1uq1"",Bjpi"B,"p"i4
RRRRRRRR)qj Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRq j)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRq 4)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR4Rq)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR)q4 )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR)Aj Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRARRjt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRRjRA)_ t)  1aRR:#H0sM:oR=)R" a1 jR";-)-" a1 jR","1)  "a4
R
RRRRRR4RA)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRA 4)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRARR4t) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRqRRBmBpqQ7_)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRqpBBm_q7Qt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRRBRqBqpm7)_Q )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR7q71jzA_ Q)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR7Rq7A1zj)_Q Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRq177z_AjQt) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRqRR7z71AQ4_)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRq177z_A4Qt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR7Rq7A1z4)_Q )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR u)tBj_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"RR-RR-Dlk0bjRHDbCHRMCsHCo#s0C
RRRRRRRR u)tBj_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRut) j _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRut) 4p_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"RRRR-R-l0kD4HRbbHCDMsCRC#oH0
CsRRRRRRRRut) 4 _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRuRR)4 t_1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRwRRA)_u :tRR0LHRR:=';j'RR--',j'"uAYq"11;''4,h" q Ap"RRRR-RR-CVC8OLN	ORNOHRbbHCDMsCRC#oH0,Cs#CNlR	OD//OCsCC#0#RNR m)tR

RRRRRqRRBmBpqu7_)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRqpBBm_q7ut) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRRBRqBqpm7)_u )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR7q71jzA_ u)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR7Rq7A1zj)_u Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRq177z_Ajut) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRqRR7z71Au4_)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRq177z_A4ut) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR7Rq7A1z4)_u )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR m)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR)Rm Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRmt) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRvRRz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"-;-Rh1YB1,qY
hBRRRRRRRRu_) p7mqRH:RMo0CC:sR=;Rj
RRRRRRRR1BqQh_ R#:R0MsHo=R:Rq"wp"1 -w-"q p1"8:RHL#NDOCRN5#HjR2;"za) C":MDNLCNRO#OH5N2#H
;S2
RRRRb
SFRs05S
SqAj,jRR:H#MR0D8_FOoH_OPC05Fs484RF0IMF2Rj;S
SqA4,4RR:H#MR0D8_FOoH_OPC05Fs484RF0IMF2Rj;S
SBQq1RH:RM0R#8F_Do_HOP0COF6s56FR8IFM0R;j2
qSSBmBpq:7RRRHM#_08DHFoOS;
S7q71RzA:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SRB :MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SiBpRH:RM0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;S S)1R a:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
Sz7maRR:FRk0#_08DHFoOC_POs0F5R668MFI0jFR2S;
S1BqmRR:FRk0#_08DHFoOC_POs0F5R668MFI0jFR22
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu7164n_..X41Rzv:FRBlMbFCRM0H0#Rs;kC
-
--------------------------1-7u_6n.4(XU---------------------------------------
vBmu mhh7aR1nu6_X.(4RU
RoRRCsMCH
O5S)Sq Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRqRR)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR q)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRAt) _iBpR#:R0MsHo=R:RY"Au1q1"-;R-AR"Y1uq1"",Bjpi"B,"p"i4
RRRRRRRR A)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRARR)_ t)  1aRR:#H0sM:oR=)R" a1 jR";-)-" a1 jR","1)  "a4
R
RRRRRR)RB Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRBRR)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR B)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRqpBBm_q7Qt) _iBpR#:R0MsHo=R:RY"Au1q1"-;R-AR"Y1uq1"",Bjpi"B,"p"i4
RRRRRRRRBqBp7mq_ Q)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRqRRBmBpqQ7_)_ t)  1aRR:#H0sM:oR=)R" a1 jR";-)-" a1 jR","1)  "a4
R
RRRRRR7Rq7A1z_ Q)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR7Rq7A1z_ Q)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRqRR7z71A)_Q )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR u)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"RR
RRRRRuRR)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR u)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRwuA_)R t:HRL0=R:R''j;-R-R''j,Y"Au1q1"4;'' ,"hpqA R"RRRRR-C-VCN8LON	RObORHDbCHRMCsHCo#s0C,l#NCDRO	C/O/#sCCN0R#)Rm Rt
RRRRR1RRmuq_)R t:HRL0=R:R''j;'--j"',AqYu1;1"',4'"q hA"p RRRRR-RR-N#FRbbHCMDHCCRso0H#C#s,NRlCO/D	OsC/C0#CRRN#qt) 
R
RRRRRRBRqBqpm7)_u Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRqRRBmBpqu7_)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRRBqBp7mq_ u)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRq177zuA_)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRq177zuA_)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR7q71_zAut) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRmRR)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRmt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR)Rm )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1h;B"-1-RY,hBqh1YBR
RRRRRR)Ru m_pq:7RR0HMCsoCRR:=jR;
RRRRRBRRq_1Q :hRRs#0HRMo:"=Rw1qp -";-q"wp"1 :HR8#DNLCNRO#jH52";Ra )z"M:CNCLDR#ONHN5O#
H2RRRRRRRRu7q7_R h:0R#soHMRR:="pwq1; "-a-")"z ,q"wp"1 
RRRRRRRR7uq77_q7A1zRL:RH:0R=jR'''--jR':N;88R''4:kR#L2
S;R
RRSR
b0FsRS5
S1q,Q:qRRRHM#_08DHFoOC_POs0F5R.n8MFI0jFR2S;
S:ARRRHM#_08DHFoOC_POs0F5R4(8MFI0jFR2S;
S:BRRRHM#_08DHFoOC_POs0F5R.68MFI0jFR2S;
S1BqQRR:H#MR0D8_FOoH_OPC05Fs686RF0IMF2Rj;S
SqpBBmRq7:MRHR8#0_oDFH
O;S7Sq7A1z,1Rq :pRRRHM#_08DHFoOS;
SRB :MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SiBpRH:RM0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;S S)1R a:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
Sz7maRR:FRk0#_08DHFoOC_POs0F5R668MFI0jFR2S;
Sq1mRF:Rk#0R0D8_FOoH_OPC05Fs.8nRF0IMF2Rj;S
SBmq1RF:Rk#0R0D8_FOoH_OPC05Fs686RF0IMF2Rj
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV761un(_.XR4U:FRBlMbFCRM0H0#Rs;kC
-
--------------------------1-7u_6n44.X.---------------------------------------
vBmu mhh7aR1nu6_X4.4R.
RoRRCsMCH
O5S)Sq Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRqRR)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR q)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRAt) _iBpR#:R0MsHo=R:RY"Au1q1"-;R-AR"Y1uq1"",Bjpi"B,"p"i4
RRRRRRRR A)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRARR)_ t)  1aRR:#H0sM:oR=)R" a1 jR";-)-" a1 jR","1)  "a4
R
RRRRRR)Ru Bt_p:iRRs#0HRMo:"=RAqYu1;1"RR--"uAYq"11,p"Bi,j""iBp4R"
RRRRRuRR)_ tB: RRs#0HRMo:"=RB" j;-R-R "Bj"",B" 4
RRRRRRRR u)t _)1R a:0R#soHMRR:="1)  "aj;-R-"1)  "aj,)R" a1 4
"
RRRRRRRRmt) _iBpR#:R0MsHo=R:RY"Au1q1"-;R-AR"Y1uq1"",Bjpi"B,"p"i4
RRRRRRRR m)t _BR#:R0MsHo=R:R "BjR";-"-RB" j, "B4R"
RRRRRmRR)_ t)  1aRR:#H0sM:oR=)R" a1 jR";-)-" a1 jR","1)  "a4
R
RRRRRRzRvp)a_ a1 _7vm RR:#H0sM:oR=1R"Y"hB-1-RY,hBqh1YB2
S;R
RRSR
b0FsRS5
S:qRRRHM#_08DHFoOC_POs0F5R448MFI0jFR2S;
S:ARRRHM#_08DHFoOC_POs0F5R448MFI0jFR2S;
SRB :MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
SiBpRH:RM0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;S S)1R a:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
Sz7maRR:FRk0#_08DHFoOC_POs0F5R.d8MFI0jFR22
S;M
C8mRBvhum ;ha
0SN0LsHkR0C#_$MLODN	F_LGVRFRu7164n_..X4RB:RFFlbM0CMRRH#0Csk;-

-------------------------7--1nu6_X.(d-n--------------------------------------m
Bvhum Rha761un(_.X
dnRRRRoCCMs5HO
qSS)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRqt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR)Rq )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR A)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR)RA Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRAt) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRBRR)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRBt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR)RB )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRR u)tp_BiRR:#H0sM:oR=AR"Y1uq1R";-"-RAqYu1,1""iBpj"",B4pi"R
RRRRRR)Ru Bt_ RR:#H0sM:oR=BR" ;j"RR--"jB "B," 
4"RRRRRRRRut) _1)  :aRRs#0HRMo:"=R)  1a;j"R"--)  1a,j"R ")14 a"R

RRRRRmRR)_ tBRpi:0R#soHMRR:="uAYq"11;-R-RY"Au1q1"B,"p"ij,p"Bi
4"RRRRRRRRmt) _RB :0R#soHMRR:="jB "-;R-BR" ,j""4B "R
RRRRRR)Rm )t_ a1 R#:R0MsHo=R:R ")1j a"-;R- ")1j a"",R)  1a
4"
RRRRRRRRpvza _)1_ av m7R#:R0MsHo=R:RY"1h;B"-1-RY,hBqh1YBR
RRRRRRqRu7 7_hRR:1Qa)h:tR=wR"q p1"-;R-)"az, ""pwq1
 "RRRRRRRRu7q7_7q71RzA:HRL0=R:R''jR'--jR':N;88R''4:kR#L;
2
b
SFRs05S
SqRR:H#MR0D8_FOoH_OPC05Fs.8nRF0IMF2Rj;S
SARR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj;S
SBRR:H#MR0D8_FOoH_OPC05Fs.86RF0IMF2Rj;S
SB: RRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;S
SBRpi:MRHR8#0_oDFHPO_CFO0sR548MFI0jFR2S;
S1)  :aRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fsn8.RF0IMF2Rj
;S2
8CMRvBmu mhh
a;S0N0skHL0#CR$LM_D	NO_GLFRRFV761un(_.XRdn:FRBlMbFCRM0H0#Rs;kC




RRRRM
C8FROlMbFC#M0;RRRRR
RR
R

