@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)qa_pYWq1
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
`

HCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0M`C
CHM8V/R/m_epQahQ_tv1
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 ap_qW1qY_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RCR0#C0_G;bs
CRRMs8bFsbC0
$

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RbbsFC$s0R1q1 _)aqqpWYX1_Zh_m_1a aX_ uu)_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5HM#k	IMFMC50#C0_G2bs2
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRR_Rqq 11)qa_pYWq1:_uR#N#CRs0bbsFC$s0R15q1a )_Wqpq_Y1uR2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHw#Rq p1"
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)qa_pYWq1Z_X__mhaa 1_u X):_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_Wqpq_Y1XmZ_h _a1 a_X_u)uR2
RRRRRCRRDR#CF_PDCFsss5_0"#0C0G_CbOsRFNM0HRM#XsRFR2Z";R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRv1_q1a )_Wqpq_Y1uN:R#l#kCsRbFsbC05$Rq 11)qa_pYWq12_u;`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )_Wqpq_Y1XmZ_h _a1 a_X_u)uR:
RRRRRNRR#l#kCsRbFsbC05$Rq 11)qa_pYWq1Z_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHM;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m




