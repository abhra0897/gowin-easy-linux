@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Wa_Qzh_hqB]h"t ;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"
`8HVCmVReQp_h_Qav
1tRRRRH0MHH
NDRRRRRPRFDM_HHl0_#0o_;/R/RDBNDER0C#RzC7sRCMVHCQ8RMRH0v#C#NRoC)0FkH
MC`8CMH/VR/pme_QQha1_vt`

HCV8VeRmp]_1q7) _7Bm R

RosCRMIH8RFI=;Rj
R
RNNDI$@#R@bR5F8#CoOCRDR	2LHCoMR
RRVRHRm5`e)p_ a1 _t1QhRqp!4=R'2LjRoLCHRM
RRRRRRHV5H!IMI8FRR&&#s0N0P_CCRM0=4=R'2L4
RRRRRRRRMIH8RFI<4=R';L4
RRRRCRRDR#CH5VRI8HMF&IR&MRC8P_CCRM0=4=R'2L4
RRRRRRRRMIH8RFI<4=R';Lj
RRRR8CM
RRRR#CDCCRLo
HMRRRRRHRIMI8FRR<=4j'L;R
RRMRC8R
RC
M8
M`C8RHV/m/Re1p_] q)7m_B7
 
`8HVCmVReqp_1)1 ah_m

RRRsRbFsbC0q$R1)1 aQ_Whh_zBh]qtu _;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5N#0sC0_P0CMRR&&!MIH82FIR4yyR55!C_M8CMPC0&R&R0f#NCLD5#0C0G_Cb2s224r*:Rf9|R->fN#0L5DC00C#_bCGs
2;RMRC8Fbsb0Cs$
R
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
bRRsCFbsR0$q 11)Wa_Qzh_hqB]h_t XmZ_ha_1q_)a he a;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
!RR5MIH82FIR>|-R55!fkH#MF	MI#M500Ns_CCPM2022R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aW_Qhz]hBq ht__XZmah_ _1a )Xu_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RIR5HFM8I|R|RN#0sC0_P0CM2-R|>!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Wa_Qzh_hqB]h_t XmZ_hh_ 7e_  _hauR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RH5IMI8F2-R|>!R55#fHkMM	F5IMC_M8CMPC0222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )_hWQ_Bzh]tqh :_uR#N#CRs0bbsFC$s0R15q1a )_hWQ_Bzh]tqh 2_u
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMERN#OMENoRC8PkNDCCRLVCFsRC0ERCCPMI0RHFM8IDROF##C"
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)Wa_Qzh_hqB]h_t XmZ_ha_1q_)a he a:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)Wa_Qzh_hqB]h_t XmZ_ha_1q_)a he a2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N#0sC0_P0CMRMOF0MNH#RRXFZsR"
2;RRRRRRRRq1_q1a )_hWQ_Bzh]tqh Z_X__mhaa 1_u X):_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)Wa_Qzh_hqB]h_t XmZ_h _a1 a_X_u)uR2
RRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RRRRRRRRq1_q1a )_hWQ_Bzh]tqh Z_X__mh _h7 he a:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)Wa_Qzh_hqB]h_t XmZ_hh_ 7e_  _hauR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0C5"MC8_P0CMRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 aQ_Whh_zBh]qtu _:#RN#CklRFbsb0Cs$qR51)1 aQ_Whh_zBh]qtu _2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqv_1)1 aQ_Whh_zBh]qtX _Zh_m_q1a) a_ea h_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 aQ_Whh_zBh]qtX _Zh_m_q1a) a_ea h_;u2
RRRRRRRRqv_1)1 aQ_Whh_zBh]qtX _Zh_m_1a aX_ uu)_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aW_Qhz]hBq ht__XZmah_ _1a )Xu_;u2
RRRRRRRRqv_1)1 aQ_Whh_zBh]qtX _Zh_m_7 h_  ehua_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aW_Qhz]hBq ht__XZm h_h 7_ea h_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_ho

CsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_CsI8HMFFI_b:CM
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRRRRRN#0sC0_P0CMRR&&!MIH82FIRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8_FIFMbCRPOFC8sC"
2;
RRRRORRFsPC_MIH8:FI
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52R`pme_1)  1a_Qqthp=R!RL4'j02REksFokEF0R
RRRRRRRRRRRRRRRRRR5RR5N#0sC0_P0CMRR&&!MIH82FIR4yy
RRRRRRRRRRRRRRRRRRRR!R5C_M8CMPC0&R&RMIH82FIRjr*:Rf9y
y4RRRRRRRRRRRRRRRRRRRRRM5C8P_CCRM0&I&RHFM8IR222R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05I8HMFOIRFsPCC28";R
RRCRRM/8R/#LNHOORFsPCN
oCRRRRC
M8
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m




