@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)a7a pq
";
V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
`8HVCmVReqp_1)1 ah_m
R
RbbsFC$s0R1q1 _)a7a pq;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RR!0f#NCLD5#0C0G_CbRs2&f&Rb0N#5e`mp _)1_ a1hQtq2p2R>|-R555545{',Ljf#bN0C50#C0_G2bs}RR-{L4'jC,0#C0_G}bs2RR&5'{4L{j,I0H8E'{4L}4}}R22>l=RHRM2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5{554j'L,Nfb#005C_#0CsGb2-}RR'{4L0j,C_#0CsGb}&2RR45{',Lj{8IH04E{'}L4}2}2RR<=l2NG
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR|2R|R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5R5545{',Lj00C#_bCGs-}RR'{4Lfj,b0N#5#0C0G_Cb}s22RR&5'{4L{j,I0H8E'{4L}4}}R22>l=RHRM2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5{554j'L,#0C0G_CbRs}-4R{',Ljf#bN0C50#C0_G2bs}&2RR45{',Lj{8IH04E{'}L4}2}2RR<=l2NG
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR;R2
CRRMs8bFsbC0
$

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RbbsFC$s0R1q1 _)a7a pqZ_X__mhaa 1_u X);_u
@RR@bR5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R555!fkH#MF	MI0M5C_#0CsGb2222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )_p7 auq_:R
RRRRRR#RN#0CsRFbsb0Cs$qR51)1 a _7p_aquC2RDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRNOEM8oCRRL$NCR8DR0NPkNDCFRM0MRHRC0ERMsNo#CRbHCOV8HCRRL$lRHMNRM8l"NG2
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)7a_ qpa__XZmah_ _1a )Xu_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)a7a pqZ_X__mhaa 1_u X)2_u
RRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R

RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRR_Rvq 11)7a_ qpa_Ru:Nk##lbCRsCFbsR0$51q1 _)a7a pq2_u;
R
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqv_1)1 a _7p_aqXmZ_h _a1 a_X_u)uR:
RRRRRNRR#l#kCsRbFsbC05$Rq 11)7a_ qpa__XZmah_ _1a )Xu_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
R`RRm_epQmth): RRoLCH:MRRDFP_MHoF
sCRRRRRRRR/8/RFFRM0MEHoR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h


`8HVCmVReBp_m)e _
mh
oRRCsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_Cs00C#_bCGsE_ONCMo:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR!0f#NCLD5#0C0G_CbRs22R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbOs_EoNMCFROPCCs8;"2
RRRRMRC8R

RRRRH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR

RRRRRPOFC0s_C_#0CsGb_D8C0NN_0H_lMR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&bRfN5#0`pme_1)  1a_Qqthp&2R&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#!f0DNLCC50#C0_G2bsR
&&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RR5{554j'L,Nfb#005C_#0CsGb2-}RR'{4L0j,C_#0CsGb}&2RR45{',Lj{8IH04E{'}L4}2}2RR==l2HMR
||RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5{554j'L,#0C0G_CbRs}-4R{',Ljf#bN0C50#C0_G2bs}&2RR45{',Lj{8IH04E{'}L4}2}2RR==l2HM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2RR
RRRRRRRRRRRRRRRRRRRR
R2RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5C"0#C0_G_bs80CDN0_N_MlHRPOFC8sC"
2;
RRRRORRFsPC_#0C0G_Cb8s_CND0__N0l:NG
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjRR&&f#bN0m5`e)p_ a1 _t1Qh2qpR
&&RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR!RRfN#0L5DC00C#_bCGs&2R&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5555'{4Lfj,b0N#5#0C0G_Cb}s2R{-R4j'L,#0C0G_Cb2s}R5&R{L4'jI,{HE80{L4'4}}}2=2R=NRlG|2R|R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5R55'{4L0j,C_#0CsGb}RR-{L4'jb,fN5#000C#_bCGs22}R5&R{L4'jI,{HE80{L4'4}}}2=2R=NRlGR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
R2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2
RRRRRRRRRRRRRRRRRRRR2R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsC_8D_0NNl0_NOGRFsPCC28";R
RRCRRMR8
RCRRM
8
RMRC8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



