@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Ba_]tqh 
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
HRRMHH0NLDRCMoH
RRRRRHV55~5NHO0FFM_MC_MI0_#NRs0=`=Rm_epQmth)h _ 1W_aaq)2|R|
RRRRRRRR5RRNHO0FFM_MC_MI0_#NRs0=`=Rm_ep)  1ah_m_Wh _q1a)Ra2|R|
RRRRRRRRRO5N0MHF__FMM_CI#s0N0=R=Re`mp)_ )_m)mhh_ 1W_aaq)2R22LHCoMR
RRRRRF_PDCFsss5_0"DQDCDoNRDPNk#CRCV0RFbsRNlsNCs0CR0NOH_FMFMM_C#I_00Ns"
2;RRRRC
M8RMRC8`

HCV8VeRmp]_1q7) _7Bm R

RosCRMIH8RFI=;Rj
HRRMo0CCHsRRj=R;R

RINDNR$#@5@RbCF#8RoCO2D	RoLCHRM
RHRRV`R5m_ep)  1aQ_1tphqRR!=4j'L2CRLo
HMRRRRRVRHRI5!HFM8I&R&RN#0sC0_P0CMRR==44'L2CRLo
HMRRRRRRRRI8HMF<IR='R4L
4;RRRRRRRRH=R<RlMk_#O	;R
RRRRRC
M8RRRRRDRC#HCRVIR5HFM8IL2RCMoH
RRRRRRRRRHV5=HR=RR4&5&RNHO0FFM_MC_MI0_#NRs0!`=Rm_ep)  1ah_m_Wh _q1a)|aR|0R#N_s0CMPC0=R!RL4'4
22RRRRRRRRRHRIMI8FRR<=4j'L;R

RRRRRHRRVNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqa&R&RN#0sC0_P0CMRR==44'L2R
RRRRRRRRRH=R<RlMk_#O	;R
RRRRRRDRC#HCRVHR5RR!=4R2
RRRRRRRRR<HR=RRH-;R4
RRRRCRRM/8R/VRHRH5IMI8F2R
RRMRC8R
RRDRC#LCRCMoH
RRRRIRRHFM8I=R<RL4'jR;
RRRRR<HR=;Rj
RRRR8CM
CRRM
8
`8CMH/VR/eRmp]_1q7) _7Bm `

HCV8VeRmp1_q1a )_
mh
bRRsCFbsR0$q 11)Ba_]tqh ;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RR#s0N0P_CCRM0&!&RI8HMFRI2|R->5ryy4k:Ml	_O#!9RfN#0L5DC00C#_bCGs;22
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 a]_Bq ht_1)  ma_ha_1q_)auR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R05#N_s0CMPC0|2R=5>R44'LRjr*:lMk_#O	-R49y
y4RRRRRRRRRRRRRRRRRRRRRf5!#L0ND0C5C_#0CsGb2|R|RN#0sC0_P0CM2
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_qB]h_t  _))m1h_aaq)_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RHRIMI8FR>|-R0!#N_s0CMPC0R;
R8CMbbsFC$s0
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRsRbFsbC0q$R1)1 a]_Bq ht__XZm1h_aaq)_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R!I8HMFRI2|R->5f!5HM#k	IMFM05#N_s0CMPC0222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Ba_]tqh Z_X__mhh_ W1)aqa;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRI8HMFRI2|R->5f!5HM#k	IMFM05#N_s0CMPC0222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Ba_]tqh Z_X__mhaa 1_u X);_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRI8HMF|IR|0R#N_s0CMPC0|2R-5>R!H5f#	kMMMFI5#0C0G_Cb2s22R;
R8CMbbsFC$s0
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
oRRCsMCN
0C
RRRR#ONCbR5sCFbs_0$0C$b2R
RRRRR`pme_1q1 R)a:CRLoRHM:PRFD#_N#0Cs
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR!=`pme_1)  ma_h _hWa_1q2)a
RRRRRRRRqRR_1q1 _)aBh]qtu _:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aBh]qtu _2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HMHR88FRM0ERONCMoRDPNkICRHH0EMkRMl	_O#$ROO#DCR0NVC#sR00NsRCCPM20";R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2R
RRRRRRRRRq1_q1a )_qB]h_t )  1ah_m_q1a)ua_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aBh]qt) _ a1 __mh1)aqa2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N10sC0RP0CMRNCPD0kNCa8R)Rz LFCVs0CRCR#0CsGbCH##FOMREoNMC28";R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp)_ )_m)mhh_ 1W_aaq)2R
RRRRRRRRRq1_q1a )_qB]h_t  _))m1h_aaq)_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a]_Bq ht_) )__mh1)aqa2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"DQDCDoNR-sCFkOOsONMCVRFRN#0sC0RP0CM"
2;
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRRRRR_Rqq 11)Ba_]tqh Z_X__mh1)aqa:_u
RRRRRRRRRRRNC##sb0RsCFbsR0$51q1 _)aBh]qtX _Zh_m_q1a)ua_2R
RRRRRRRRRR#CDCPRFDs_Cs_Fs0#5"00Ns_CCPMO0RFNM0HRM#XsRFR2Z";R
RRRRRRHRRVNR5OF0HMM_F_IMC_N#0s!0R=mR`eQp_t)hm  _hWa_1q2)a
RRRRRRRRRRRq1_q1a )_qB]h_t XmZ_h _hWa_1q_)auR:
RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a]_Bq ht__XZmhh_ 1W_aaq)_
u2RRRRRRRRRCRRDR#CF_PDCFsss5_0"N#0sC0_P0CMRMOF0MNH#RRXFZsR"
2;RRRRRRRRRqq_1)1 a]_Bq ht__XZmah_ _1a )Xu_
u:RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_qB]h_t XmZ_h _a1 a_X_u)uR2
RRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_ep)  1ah_m_Wh _q1a)
a2RRRRRRRRR_Rvq 11)Ba_]tqh :_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)Ba_]tqh 2_u;R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2R
RRRRRRRRRv1_q1a )_qB]h_t )  1ah_m_q1a)ua_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aBh]qt) _ a1 __mh1)aqa2_u;R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp)_ )_m)mhh_ 1W_aaq)2R
RRRRRRRRRv1_q1a )_qB]h_t  _))m1h_aaq)_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a]_Bq ht_) )__mh1)aqa2_u;


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRRRRv1_q1a )_qB]h_t XmZ_ha_1q_)auR:
RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a]_Bq ht__XZm1h_aaq)_;u2
RRRRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R!Re`mpt_Qh m)_Wh _q1a)
a2RRRRRRRRRvRR_1q1 _)aBh]qtX _Zh_m_Wh _q1a)ua_:R
RRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qB]h_t XmZ_h _hWa_1q_)au
2;RRRRRRRRRvRR_1q1 _)aBh]qtX _Zh_m_1a aX_ uu)_:R
RRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qB]h_t XmZ_h _a1 a_X_u)u
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
V`H8RCVm_epB me)h_m
C
oMNCs0
C
RRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR

RRHV5pme_eBm A)_qB1Q_2mhRoLCH:MRRDFP_POFCLs_NO#H
R
RRFROP_CsI8HMFFI_b:CM
RRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&RR
RRRRRRRRRRRRRRRRR0R#N_s0CMPC0&R&RH!IMI8F2
R2RRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05I8HMFFI_bRCMOCFPs"C82R;
R
RRRRRROCFPsH_IMI8F_FOD#
C:RRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRI8HMF&IR&HR5RR==4&R&RO5N0MHF__FMM_CI#s0N0=R!Re`mp _)1_ amhh_ 1W_aaq)RR||#s0N0P_CCRM0!4=R'2L4222R
RRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8_FIO#DFCFROPCCs8;"2
CRRM/8R/#LNHOORFsPCN
oC
RRRH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR

RHRRVNR5OF0HMM_F_IMC_N#0s=0R=mR`e)p_ a1 __mhh_ W1)aqaL2RCMoHRF:RPOD_FsPC_MIH8_FIsCC#0R#
RRRRRPOFCIs_HFM8IC_s##C0:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRR0R#N_s0CMPC0&R&RMIH82FIRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8_FIsCC#0O#RFsPCC28";R
RRMRC8R
RR8CMRO//FCsMsFROPNCso
CR
MRC8/R/Rpme_eBm h)_m
h 
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m
