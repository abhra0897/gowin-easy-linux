@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)awv)q 
";
V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
RMRHHN0HDCRLo
HMRRRRH5VR~N55OF0HMM_F_IMC_N#0s=0R=mR`eQp_t)hm  _hWa_1q2)aR
||RRRRRRRRRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2|R|
RRRRRRRRNR5OF0HMM_F_IMC_N#0s=0R=mR`e p_)))m__mhh_ W1)aqa222RoLCHRM
RRRRRPRFDs_Cs_Fs0Q5"DoDCNPDRNCDkR0#CRsVFRsbNN0lCCNsROF0HMM_F_IMC_N#0s20";R
RRMRC8R
RRVRHRN5lG	_O#&R&RN5lG	_O#RR<l_HMO2	#2CRLo
HMRRRRRFRRPCD_sssF_"05QCDDoRNDbNNslCC0sNRPD#kCR0#CRCIEslCRHOM_	>#RRGlN_#O	"
2;RRRRC
M8RMRC8`

HCV8VeRmp1_q1a )_
mh
HRRMo0CCHsRHRR=jR;
RosCRMIHRj=R;R
RsRCos0_#N_s0CMPC0RR=j
;
RDRNI#N$R5@@bCF#8RoCO2D	RoLCHRM
RsRR_N#0sC0_P0CMRR<=#s0N0P_CC;M0
CRRM
8
RDRNI#N$R5@@bCF#8RoCO2D	RoLCHRM
RHRRV`R5m_ep)  1aQ_1tphqRR!=44'L2CRLo
HMRRRRRHRHRR<=jR;
RRRRRMIHRR<=jR;
RCRRMR8
RCRRDR#CLHCoMR
RRRRRH5VRl_NGOR	#>2RjRoLCHRM
RRRRRORRNR#C5MIH2RR
RRRRRRRRRRj:LHCoMR
RRRRRRRRRRVRHR_5s#s0N0P_CCRM0=4=R'RLj&#&R00Ns_CCPM=0R='R4L&4R&R
RRRRRRRRRRRRRR0R5C_#0CsGbRR!=44'L2L2RCMoH
RRRRRRRRRRRRIRRH<MR='R4L
4;RRRRRRRRRRRRRHRHRR<=l_NGO;	#
RRRRRRRRRRRR8CM
RRRRRRRRCRRMR8
RRRRRRRRRR4:LHCoMR
RRRRRRRRRRVRHR_5s#s0N0P_CCRM0=4=R'RLj&#&R00Ns_CCPM=0R='R4L&4R&R
RRRRRRRRRRRRRRORN0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)R
&&RRRRRRRRRRRRRRRR00C#_bCGs=R!RL4'4L2RCMoH
RRRRRRRRRRRRHRRH=R<RGlN_#O	;R
RRRRRRRRRRMRC8R
RRRRRRRRRRDRC#HCRVHR5H=R<R|4R|CR0#C0_GRbs=4=R'2L4RoLCHRM
RRRRRRRRRRRRRMIHRR<=4j'L;R
RRRRRRRRRRMRC8R
RRRRRRRRRRDRC#LCRCMoH
RRRRRRRRRRRRHRRH=R<RRHH-
4;RRRRRRRRRRRRC
M8RRRRRRRRRMRC8R
RRRRRRMRC8#ONCR
RRRRRC
M8RRRRRDRC#HCRVlR5HOM_	>#RRRj2LHCoMR
RRRRRRNRO#5CRI2HMRR
RRRRRRRRRjL:RCMoH
RRRRRRRRRRRRRHV5#s_00Ns_CCPM=0R='R4L&jR&0R#N_s0CMPC0=R=RL4'4&R&
RRRRRRRRRRRRRRRRC50#C0_GRbs!4=R'2L42CRLo
HMRRRRRRRRRRRRRHRIM=R<RL4'4R;
RRRRRRRRRRRRRRHH<l=RHOM_	
#;RRRRRRRRRRRRC
M8RRRRRRRRRMRC8R
RRRRRRRRR4L:RCMoH
RRRRRRRRRRRRRHV5#s_00Ns_CCPM=0R='R4L&jR&0R#N_s0CMPC0=R=RL4'4&R&RR
RRRRRRRRRRRRRRORN0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)R
&&RRRRRRRRRRRRRRRR00C#_bCGs=R!RL4'4L2RCMoH
RRRRRRRRRRRRHRRH=R<RMlH_#O	;R
RRRRRRRRRRMRC8R
RRRRRRRRRRDRC#HCRVHR5H=R<R|4R|CR0#C0_GRbs=4=R'2L4RoLCHRM
RRRRRRRRRRRRRMIHRR<=4j'L;R
RRRRRRRRRRMRC8R
RRRRRRRRRRDRC#LCRCMoH
RRRRRRRRRRRRHRRH=R<RRHH-
4;RRRRRRRRRRRRC
M8RRRRRRRRRMRC8R
RRRRRRMRC8#ONCR
RRRRRC
M8RRRRC
M8RMRC8R

RFbsb0Cs$1Rq1a )_qw)vv _Q_hjvjqX_
u;R@R@5#bFCC8oR	OD2RR
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
fRRsCF#5N#0sC0_P0CM2-R|>CR0#C0_G;bs
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 a)_wq_v  _))m1h_aaq)_
u;R@R@5#bFCC8oR	OD2RR
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
!RR5Ffs##C500Ns_CCPMR02&I&RH;M2
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 a)_wq_v v_QhBB] i;_u
@RR@F5b#oC8CDRO	
2RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5Ffs##C500Ns_CCPMR02&!&RI2HMR>|-R!5500C#_bCGslr*HOM_	2#92R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)awv)q q_vX]_B _BiuR;
R5@@bCF#8RoCO2D	RR
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RfR5sCF#5N#0sC0_P0CM2&R&RH!IM|2R-5>R!#0C0G_Cb*srjN:lG	_O#y9Ry04RC_#0CsGb2R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)awv)q  _)1_ am1h_aaq)_hvQ_ B]Bui_;R
R@b@5F8#CoOCRDR	2
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RFfs##C500Ns_CCPMR02|R->5C!0#C0_GRbsy
y4RRRRRRRRRRRRRRRRRRRRRRRRR5R5!#0C0G_Cb*sr5MlH_#O	Rj>RRl?RHOM_	4#-R4:R2R92FRs
RRRRRRRRRRRRRRRRRRRRRRRRR!R500C#_bCGsjr*:H5lM	_O#RR>jRR?l_HMO-	#4RR:4R29yRyjf#sFC05#N_s0CMPC0222
RRRRRRRRRRRRRRRRRRRRRRRR;R2
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 a)_wq_v )  1ah_m_q1a)va_qBX_]i B_
u;R@R@5#bFCC8oR	OD2RR
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRf#sFC05#N_s0CMPC0&2R&0R!C_#0CsGb2=R|>!R500C#_bCGsjr*:N5lG	_O#RR>jRR?l_NGO-	#4RR:4R29y
y4RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0R5C_#0CsGbRR||5Ffs##C500Ns_CCPM2022R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2RR;R
RCbM8sCFbs
0$
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRsRbFsbC0q$R1)1 a)_wq_v XmZ_ha_1q_)auR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R!RR5MIH2-R|>!R55#fHkMM	F5IM#s0N0P_CC2M02
2;RRRRCbM8sCFbs
0$
RRRRFbsb0Cs$1Rq1a )_qw)vX _Zh_m_Wh _q1a)ua_;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RRIR5HRM2|R->5f!5HM#k	IMFM05#N_s0CMPC0222;R
RRMRC8Fbsb0Cs$R

RbRRsCFbsR0$q 11)wa_) qv__XZmah_ _1a )Xu_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5RR5f#sFC05#N_s0CMPC0&2&5H!IM22RRR||5MIH2RR2|R->5f!5HM#k	IMFMC50#C0_G2bs2
2;RRRRCbM8sCFbs
0$
RRRRFbsb0Cs$1Rq1a )_qw)vv _QXh_Z]_B _BiuR;
R@RR@F5b#oC8CDRO	R2
R8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R5RRf#sFC05#N_s0CMPC0&2R&IR!HRM2|R->5!555#fHkMM	F5IM00C#_bCGs222rH*lM	_O#292;R
RRMRC8Fbsb0Cs$R

RbRRsCFbsR0$q 11)wa_) qv__XZvjQh_Xvqj;_u
RRRR5@@bCF#8RoCO2D	
RRRR#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRRFfs##C500Ns_CCPMR02|R->5f!5HM#k	IMFMC50#C0_G2bs2
2;RRRRCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRH5VRl_HMOR	#=j=RRR&&l_NGOR	#=j=R2CRLoRHM:_RNNC##sV0_sCNl_MlHjN_lGRj
RRRRRRRRRqq_1)1 a)_wq_v vjQh_Xvqj:_u
RRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_) qv_hvQjq_vXuj_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHR0MFRza) ERIHRDC#s0N0PRCCRM0HN#R#s#C0RC8IMECR0LFENRbsCNl0#CsRMlH_#O	R8NMRGlN_#O	RCNsR0#CRR0Fj;"2
RRRRRRRR8CM
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_hQtm_) h_ W1)aqa|R|
RRRRRRRRRRRR0NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)aRoLCH:MRRHN_osMFCs_F_sCsFFs_MC_MI0_#N
s0RRRRRRRRRVRHRH5lM	_O#RR>jL2RCMoHRN:R_#N#C_s0VlsNCH_lME_OC
O	RRRRRRRRRRRRq1_q1a )_qw)vv _QBh_]i B_
u:RRRRRRRRRRRRNC##sb0RsCFbsR0$51q1 _)awv)q Q_vh]_B _Biu
2RRRRRRRRRRRRRCCD#RDFP_sCsF0s_5C"a#C0RGCbs#F#HM#RHRza) CRLVCFsRNCDbR#CF#VRbHCOV8HCRMlHHllkRMlH_#O	ROO$DRC#VlsFRN#0sC0RP0CM"
2;RRRRRRRRRMRC8R
RRRRRRRRRH5VRl_NGOR	#>2RjRoLCH:MRRNN_#s#C0s_VN_lCl_NGOOEC	R
RRRRRRRRRR_Rqq 11)wa_) qv_Xvq_ B]Bui_:R
RRRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a)_wq_v v_qXBB] i2_uRR
RRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHM#RFa0R)Rz IEH0H#MRbHCOV8HCRGlNHllkRGlN_#O	ROO$DRC#VlsFRN#0sC0RP0CM"
2;RRRRRRRRRMRC8R
RRRRRRMRC8R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2CRLoRHM:_RNsCC#0M_F_IMC_N#0sR0
RRRRRRRRRRHV5MlH_#O	Rj>R2CRLoRHM:_RNNC##sV0_sCNl_#sCCF0_M0_#N_s0l_HMOOEC	R
RRRRRRRRRR_Rqq 11)wa_) qv_1)  ma_ha_1q_)av_QhBB] i:_u
RRRRRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_qw)v) _ a1 __mh1)aqaQ_vh]_B _BiuR2
RRRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRRH#a )zRVLCFRsCCbDN#FCRVbR#CVOHHRC8lHHMlRkll_HMOR	#OD$OCV#RsRFl#s0N0PRCC"M02R;
RRRRRRRRR8CM
RRRRRRRRHRRVlR5NOG_	>#RRRj2LHCoMRR:N#_N#0Cs_NVslsC_C0#C__FM#s0N0N_lGE_OC
O	RRRRRRRRRRRRq1_q1a )_qw)v) _ a1 __mh1)aqaq_vX]_B _BiuR:
RRRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_) qv_1)  ma_ha_1q_)av_qXBB] i2_u
RRRRRRRRRRRR#CDCPRFDs_Cs_Fs0a5"CR#0CsGbCH##FHMR#FRM0)RazI RHH0EMbR#CVOHHRC8lHNGlRkll_NGOR	#OD$OCV#RsRFl#s0N0PRCC"M02R;
RRRRRRRRR8CM
RRRRRRRR8CM
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)aRoLCH:MRRCN_sssF__FMM_CI#s0N0R
RRRRRRRRRq1_q1a )_qw)v  _)m)_ha_1q_)auR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_qw)v  _)m)_ha_1q_)auR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0Q5"DoDCN#DR00NsRCCPMI0REEHOR#ENRFsCOsOkCL8RCsVFCFROlCbD0MHFRRFVOsksCRM0I8HMF2I";R
RRRRRRMRC8


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 a)_wq_v XmZ_ha_1q_)auR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_) qv__XZm1h_aaq)_
u2RRRRRRRRCCD#RDFP_sCsF0s_50"#N_s0CMPC0FROMH0NMX#RRRFsZ;"2
R
RRRRRRVRHRl5RNOG_	>#RR2jRRoLCH:MRRNN_#s#C0s_VN_lCGFx_MC_0#C0_G
bsRRRRRRRRR_Rqq 11)wa_) qv__XZmah_ _1a )Xu_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a)_wq_v XmZ_h _a1 a_X_u)uR2
RRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;
RRRRRRRRHRRVNR5OF0HMM_F_IMC_N#0s!0R=mR`eQp_t)hm  _hWa_1qR)a2CRLoRHM:_RNNC##sV0_sCNl__GxFMM_C#I_00Ns
RRRRRRRRRRRRqq_1)1 a)_wq_v XmZ_h _hWa_1q_)auR:
RRRRRRRRRNRR#s#C0sRbFsbC05$Rq 11)wa_) qv__XZmhh_ 1W_aaq)_
u2RRRRRRRRRRRRCCD#RDFP_sCsF0s_50"#N_s0CMPC0FROMH0NMX#RRRFsZ;"2
RRRRRRRRCRRMR8
RRRRRCRRMR8
RRRRRCRRDR#CH5VRRMlH_#O	Rj>RRL2RCMoHRN:R_#N#C_s0VlsNCH_lMx_G_COEOR	
RRRRRRRRRqq_1)1 a)_wq_v v_QhXBZ_]i B_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 a)_wq_v v_QhXBZ_]i B_
u2RRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
R
RRRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_epQmth)h _ 1W_aaq)RL2RCMoHRN:R_#N#C_s0VlsNCx_G__FMM_CI#s0N0R
RRRRRRRRRR_Rqq 11)wa_) qv__XZmhh_ 1W_aaq)_
u:RRRRRRRRRRRRNC##sb0RsCFbsR0$51q1 _)awv)q Z_X__mhh_ W1)aqa2_u
RRRRRRRRRRRR#CDCPRFDs_Cs_Fs0#5"00Ns_CCPMO0RFNM0HRM#XsRFR2Z";R
RRRRRRRRRC
M8RRRRRRRRC
M8RRRRRRRRCCD#RoLCH:MRRNN_#s#C0s_VN_lCGlx_H_MjljNGRR//5lR5HOM_	=#R=2RjRR&&5GlN_#O	RR==j22R
RRRRRRRRqRR_1q1 _)awv)q Z_X_hvQjq_vXuj_:R
RRRRRRRRRNC##sb0RsCFbsR0$51q1 _)awv)q Z_X_hvQjq_vXuj_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RRRRRCRRMR8
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRH5VRl_HMOR	#=j=RRR&&l_NGOR	#=j=R2CRLoRHM:_RlNC##sV0_sCNl_MlHjN_lGRj
RRRRRRRRRqv_1)1 a)_wq_v vjQh_Xvqj:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)wa_) qv_hvQjq_vXuj_2R;
RRRRRCRRMR8
RRRRRHRRVNR5OF0HMM_F_IMC_N#0s=0R=mR`eQp_t)hm  _hWa_1qR)a|R|
RRRRRRRRRNRROF0HMM_F_IMC_N#0s=0R=mR`e p_)))m__mhh_ W1)aqaL2RCMoHRl:R_MHoF_sCFCs_sssF__FMM_CI#s0N0R
RRRRRRRRRH5VRl_HMOR	#>2RjRoLCH:MRRNl_#s#C0s_VN_lCl_HMOOEC	R
RRRRRRRRRR_Rvq 11)wa_) qv_hvQ_ B]Bui_:R
RRRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a)_wq_v v_QhBB] i2_u;R
RRRRRRRRRC
M8RRRRRRRRRVRHRN5lG	_O#RR>jL2RCMoHRl:R_#N#C_s0VlsNCN_lGE_OC
O	RRRRRRRRRRRRv1_q1a )_qw)vv _qBX_]i B_
u:RRRRRRRRRRRRNk##lbCRsCFbsR0$51q1 _)awv)q q_vX]_B _Biu
2;RRRRRRRRRMRC8R
RRRRRRMRC8R
RRRRRRVRHRO5N0MHF__FMM_CI#s0N0=R=Re`mp _)1_ amhh_ 1W_aaq)2CRLoRHM:_RlsCC#0M_F_IMC_N#0sR0
RRRRRRRRRRHV5MlH_#O	Rj>R2CRLoRHM:_RlNC##sV0_sCNl_#sCCF0_M0_#N_s0l_HMOOEC	R
RRRRRRRRRR_Rvq 11)wa_) qv_1)  ma_ha_1q_)av_QhBB] i:_u
RRRRRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qw)v) _ a1 __mh1)aqaQ_vh]_B _Biu
2;RRRRRRRRRMRC8R
RRRRRRRRRH5VRl_NGOR	#>2RjRoLCH:MRRNl_#s#C0s_VN_lCsCC#0M_F_N#0sl0_NOG_EiCO
RRRRRRRRRRRRqv_1)1 a)_wq_v )  1ah_m_q1a)va_qBX_]i B_
u:RRRRRRRRRRRRNk##lbCRsCFbsR0$51q1 _)awv)q  _)1_ am1h_aaq)_Xvq_ B]Bui_2R;
RRRRRRRRR8CM
RRRRRRRR8CM
RRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR==`pme_) )mm)_h _hWa_1q2)aRoLCH:MRRCl_sssF__FMM_CI#s0N0R
RRRRRRRRRv1_q1a )_qw)v  _)m)_ha_1q_)auR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qw)v  _)m)_ha_1q_)au
2;RRRRRRRRC
M8
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRvRR_1q1 _)awv)q Z_X__mh1)aqa:_u
RRRRRRRR#N#kRlCbbsFC$s0R15q1a )_qw)vX _Zh_m_q1a)ua_2
;
RRRRRRRRH5VRRGlN_#O	Rj>RRL2RCMoHRl:R_#N#C_s0VlsNCx_G__FM00C#_bCGsR
RRRRRRRRRv1_q1a )_qw)vX _Zh_m_1a aX_ uu)_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)awv)q Z_X__mhaa 1_u X)2_u;R

RRRRRRRRRRHV50NOH_FMFMM_C#I_00NsRR!=`pme_hQtm_) h_ W1)aqaRR2LHCoMRR:l#_N#0Cs_NVslGC_xM_F_IMC_N#0sb0_
RRRRRRRRRRRRqv_1)1 a)_wq_v XmZ_h _hWa_1q_)auR:
RRRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)wa_) qv__XZmhh_ 1W_aaq)_;u2
RRRRRRRRCRRMR8
RRRRRCRRMR8
RRRRRCRRDR#CH5VRRMlH_#O	Rj>RRL2RCMoHRl:R_#N#C_s0VlsNCH_lMx_G_COEOR	
RRRRRRRRRqv_1)1 a)_wq_v v_QhXBZ_]i B_
u:RRRRRRRRR#RN#CklRFbsb0Cs$qR51)1 a)_wq_v v_QhXBZ_]i B_;u2
R
RRRRRRRRRH5VRNHO0FFM_MC_MI0_#NRs0!`=Rm_epQmth)h _ 1W_aaq)RL2RCMoHRl:R_#N#C_s0VlsNCx_G__FMM_CI#s0N0R
RRRRRRRRRR_Rvq 11)wa_) qv__XZmhh_ 1W_aaq)_
u:RRRRRRRRRRRRNk##lbCRsCFbsR0$51q1 _)awv)q Z_X__mhh_ W1)aqa2_u;R
RRRRRRRRRC
M8RRRRRRRRC
M8RRRRRRRRCCD#RoLCH:MRRNl_#s#C0s_VN_lCGlx_H_MjljNGRR//5lR5HOM_	=#R=2RjRR&&5GlN_#O	RR==j22R
RRRRRRRRvRR_1q1 _)awv)q Z_X_hvQjq_vXuj_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)awv)q Z_X_hvQjq_vXuj_2R;
RRRRRCRRMR8
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epQmth): RRoLCH:MRRDFP_MHoF
sCRRRRRRRR/8/RFFRM0MEHo
R;RRRRRMRC8R
RRRRR8NCVkRD0RRRR:MRHHN0HDPRFDs_Cs_Fs0"5"2R;
RCRRMN8O#
C
RMRC8MoCC0sNC`

CHM8V/R/Rpme_1q1 _)am
h
`8HVCmVReBp_m)e _
mh
oRRCsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _1AqQmB_hL2RCMoHRF:RPOD_FsPC_#LNH
O
RRRRRFROP_CsVlsNC0_#N:s0
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52R`pme_1)  1a_Qqthp=R!RL4'j&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RRf#sFC05#N_s0CMPC02222R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05#s0N0P_CCRM0OCFPs"C82R;
RRRRC
M8RRRRC
M8
CRRMC8oMNCs0
C
`8CMH/VR/eRmpm_Be_ )m
h

