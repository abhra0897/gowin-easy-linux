context IEEE_BIT_CONTEXT is
     library IEEE;
     use IEEE.NUMERIC_BIT.all;
end context IEEE_BIT_CONTEXT;
