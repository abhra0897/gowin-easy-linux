context IEEE_STD_CONTEXT is
     library IEEE;
     use IEEE.STD_LOGIC_1164.all;
     use IEEE.NUMERIC_STD.all;
end context IEEE_STD_CONTEXT;
