@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Wa_Qmh7W
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
V`H8RCVm_ep1)]q B7_m
7 
sRRCIoRHFM8IRR=j
;
RDRNI#N$RR@@5#bFCC8oR	OD2CRLo
HMRRRRH5VR`pme_1)  1a_Qqthp=R!RL4'jL2RCMoH
RRRRHRRV!R5I8HMF&IR&0R#N_s0CMPC0=R=RL4'4R2
RRRRRIRRHFM8I=R<RL4'4R;
RRRRR#CDCVRHRH5IMI8FRR&&C_M8CMPC0=R=RL4'4R2
RRRRRIRRHFM8I=R<RL4'jR;
RCRRMR8
RCRRDR#CLHCoMR
RRRRRI8HMF<IR='R4L
j;RRRRC
M8RMRC8`

CHM8V/R/Rpme_q1])_ 7B m7
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 aQ_WhW7m_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R#R500Ns_CCPM&0R&IR!HFM8Iy2Ry54R!M5C8P_CCRM0&0&RC_#0CsGb2*2r49:fR>|-R#0C0G_Cb
s;RMRC8Fbsb0Cs$`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRsRbFsbC0q$R1)1 aQ_WhW7m__XZm1h_aaq)_  ehua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R!H5IMI8F2-R|>!R55#fHkMM	F5IM#s0N0P_CC2M02
2;RMRC8Fbsb0Cs$R

RFbsb0Cs$1Rq1a )_hWQ7_mWXmZ_h _a1 a_X_u)uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
RH5IMI8F2-R|>!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Wa_Qmh7WZ_X__mh _h7 he a;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RRI8HMFRI2|R->5f!5HM#k	IMFMM5C8P_CC2M02
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRR_Rqq 11)Wa_Qmh7W:_uR#N#CRs0bbsFC$s0R15q1a )_hWQ7_mWuR2
RRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMOMENoRC8PkNDCkR8soHMRRNMFMbCRCCPMI0RHFM8I;"2
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)Wa_Qmh7WZ_X__mh1)aqae_  _hauR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_hWQ7_mWXmZ_ha_1q_)a he a2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N#0sC0_P0CMRMOF0MNH#RRXFZsR"
2;RRRRRRRRq1_q1a )_hWQ7_mWXmZ_h _a1 a_X_u)uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_hWQ7_mWXmZ_h _a1 a_X_u)uR2
RRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RRRRRRRRq1_q1a )_hWQ7_mWXmZ_hh_ 7e_  _hauR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_hWQ7_mWXmZ_hh_ 7e_  _hauR2
RRRRRRRRR#CDCPRFDs_Cs_Fs0C5"MC8_P0CMRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 aQ_WhW7m_Ru:Nk##lbCRsCFbsR0$51q1 _)aW7QhmuW_2
;

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rvq 11)Wa_Qmh7WZ_X__mh1)aqae_  _hauR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )_hWQ7_mWXmZ_ha_1q_)a he a2_u;R
RRRRRR_Rvq 11)Wa_Qmh7WZ_X__mhaa 1_u X):_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)Wa_Qmh7WZ_X__mhaa 1_u X)2_u;R
RRRRRR_Rvq 11)Wa_Qmh7WZ_X__mh _h7 he a:_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)Wa_Qmh7WZ_X__mh _h7 he a2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
R
RRVRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRRRH5VRm_epB me)q_A1_QBmRh2LHCoMRR:F_PDOCFPsN_L#
HO
RRRRORRFsPC_MIH8_FIFMbC:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRR0R#N_s0CMPC0&R&RH!IMI8F2
R2RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5H"IMI8F_CFbMFROPCCs8;"2
R
RRRRROCFPsH_IMI8F:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25e`mp _)1_ a1hQtq!pR='R4LRj20FEskFoEkR0
RRRRRRRRRRRRRRRRRRRR505#N_s0CMPC0&R&RH!IMI8F2yRy4R
RRRRRRRRRRRRRRRRRR5RR!8CM_CCPM&0R&HRIMI8F2*Rrj9:fR4yy
RRRRRRRRRRRRRRRRRRRRCR5MC8_P0CMRR&&I8HMF2I2RR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"MIH8RFIOCFPs"C82R;
RRRRCRM8/N/L#RHOOCFPsCNo
RRRR8CM
M
C8MoCC0sNC`

CHM8V/R/Rpme_eBm m)_h



