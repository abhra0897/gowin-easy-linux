@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11))a_q ht"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
`8HVCmVReqp_1)1 ah_m
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
RRRsRbFsbC0q$R1)1 aq_)h_t uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R55500C#_bCGs=R>RMlH2&R&RC50#C0_GRbs<l=RN2G2RR!=4j'L2R;
R8CMbbsFC$s0
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RbRRsCFbsR0$q 11))a_q ht__XZmah_ _1a )Xu_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5f!5HM#k	IMFMC50#C0_G2bs2
2;RRRRCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )_h)qtu _:#RN#0CsRFbsb0Cs$qR51)1 aq_)h_t uC2RDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRNCPD0kNC0#RFRRNPkNDCkRF08#HCER0CNRsMRoC#ObCHCVH8$RLRsbNN0lCCRs#lRHMNRM8l"NG2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRq1_q1a )_h)qtX _Zh_m_1a aX_ uu)_:RR
RRRRR#RN#0CsRFbsb0Cs$qR51)1 aq_)h_t XmZ_h _a1 a_X_u)uR2
RRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRR_Rvq 11))a_q ht_Ru:Nk##lbCRsCFbsR0$51q1 _)a)tqh 2_u;`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRRqv_1)1 aq_)h_t XmZ_h _a1 a_X_u)uR:
RRRRRRRRNk##lbCRsCFbsR0$51q1 _)a)tqh Z_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
R
RRVRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRRRH5VRm_epB me)q_1hYQa_2mhRoLCH:MRRDFP_POFC#s_N0MH$R

RRRRRPOFC0s_C_#0CsGb_NOEM:oC
RRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRRRRR#!f0DNLCC50#C0_G2bsR22R
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_NOEMRoCOCFPs"C82R;
RRRRCRM8/N/#M$H0RPOFCosNCR

RRRRH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR
R
RRRRORRFsPC_#0C0G_CbNs_0H_lMR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRRRRRRRRRRRRRRfRRsCF#5#0C0G_Cb=sR=HRlM22RRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbNs_0H_lMFROPCCs8;"2
R
RRRRROCFPsC_0#C0_G_bsNl0_N
G:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRf#sFCC50#C0_GRbs=l=RNRG22
R2RRRRRRRRRRRRRRRRRRRRRDFP_POFC0s_5C"0#C0_G_bsNl0_NOGRFsPCC28";R
RRCRRMR8
RCRRM
8
CoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
