@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11) a_e_ huQq)a;Y"
R
R`OHMDCk8R0"#8P_FDN_0#E	3"`

HCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0M`C
CHM8V/R/m_epQahQ_tv1
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 ae_  uh_qa)QY;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
5RR!55^00C#_bCGs222;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_  ehq_u)YQa__XZmah_ _1a )Xu_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R5!H5f#	kMMMFI5#0C0G_Cb2s22
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRR_Rqq 11) a_e_ huQq)auY_:#RN#0CsRFbsb0Cs$qR51)1 ae_  uh_qa)QY2_u
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCPRFDs_Cs_Fs0a5"CR#0CsGbCH##F8MRFRC#MRF0CHGELRH0CMPCRsbNH"0$2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 ae_  uh_qa)QYZ_X__mhaa 1_u X):_u
RRRRRRRR#N#CRs0bbsFC$s0R15q1a )_  ehq_u)YQa__XZmah_ _1a )Xu_
u2RRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 ae_  uh_qa)QY:_uR#N#kRlCbbsFC$s0R15q1a )_  ehq_u)YQa_;u2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRvRR_1q1 _)a he _)uqQ_aYXmZ_h _a1 a_X_u)uR:
RRRRRNRR#l#kCsRbFsbC05$Rq 11) a_e_ huQq)aXY_Zh_m_1a aX_ uu)_2R;
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epQmth): RRoLCH:MRRDFP_MHoF
sCRRRRRRRR/8/RFFRM0MEHo
R;RRRRRMRC8R
RRRRR8NCVkRD0RRRR:MRHHN0HDPRFDs_Cs_Fs0"5"2R;
RCRRMN8O#
C
RMRC8MoCC0sNC`

CHM8V/R/Rpme_1q1 _)am
h
`8HVCmVReBp_m)e _
mh
MoCC0sNCR

RHRRVOR5FsPCN_oCDCCPD=R!Re`mpm_Be_ )h mh2CRLoRHM:PRFDF_OP
CsRRRRRRHV5pme_eBm 1)_qahQYh_m2CRLoRHM:PRFDF_OP_Cs#HNM0R$

RRRRORRFsPC_#0C0G_CbOs_EoNMCR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R55R`pme_1)  1a_Qqthp=R!RL4'j&2R&R
RRRRRRRRRRRRRRRRRR!RRfN#0L5DC00C#_bCGs22RRR2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbOs_EoNMCFROPCCs8;"2
RRRRMRC8/R/#HNM0O$RFsPCN
oCRRRRC
M8
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m
