@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Za_ _)mm_h ]"ma;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"
RHR`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCR
R`8CMH
V
`8HVCmVReqp_1)1 ah_m
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RbRRsCFbsR0$q 11)Za_ _)mm_h ]_maXuZ_;R
RR@R@5#bFCC8oR	OD2R
RRHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RR!R55#fHkMM	F5IM00C#_bCGs222;R
RRMRC8Fbsb0Cs$R
R`8CMH/VR/eRmpv_QuBpQQXa_BB] iw_mwC
`MV8HRR//m_epX B]Bmi_w
w
RsRbFsbC0q$R1)1 a _Z)mm_h] _mua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R!H5f#	kMMMFI5#0C0G_Cb2s2R>|-RF5fMFCE00j5C_#0CsGb2
2;RMRC8Fbsb0Cs$R

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)aZm )_ mh_a]m_Ru:RNRR#s#C0sRbFsbC05$Rq 11)Za_ _)mm_h ]_mauR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRMOF0MNH#FRls0CRERNM4#RN#0CsCL8RH"0#2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 a _Z)mm_h] _mXa_Z:_uR#N#CRs0bbsFC$s0R15q1a )_)Z mh_m m_]aZ_X_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2R;
RM`C8RHV/m/ReQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/Rpme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRR_Rvq 11)Za_ _)mm_h ]_mauR:RR#RN#CklRFbsb0Cs$qR51)1 a _Z)mm_h] _mua_2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqv_1)1 a _Z)mm_h] _mXa_Z:_uR#N#kRlCbbsFC$s0R15q1a )_)Z mh_m m_]aZ_X_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/RR/FR7R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
RRRRRHRIsrCRI0H8E:-4j09RC_#0CsGb_=4RR#0C0G_Cb-sRRI{{HE80-44{'}Lj}',4L;4}
RRRRsRRCroRI0H8E:-4jF9RMEC_F_0#OOEC	;C8
C
oMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )1QqhamY_hL2RCMoHRF:RPOD_FsPC_M#NH
0$
RRRRORRFsPC_#0C0G_CbOs_EoNMCR:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	R`55m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRfR!#L0ND0C5C_#0CsGb22R2
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_NOEMRoCOCFPs"C82R;
RRRRCRM8/N/#M$H0RPOFCosNCR

RRRRH5VRm_epB me)m_B))h _2mhRoLCH:MRRDFP_POFCOs_FCsMsR

RRRRRINDNR$#@b@5F8#CoOCRDR	2LHCoMR
RRRRRRVRHRm5`e)p_ a1 _t1QhRqp!4=R'2LjRoLCHRM
RRRRRRRRRRHV5C50#C0_GRbs^CR0#C0_G2bs=I={HE80{L4'j2}}RoLCHRM
RRRRRRRRRHRRV5R500C#_bCGsRR&00C#_bCGs2_4RR=={8IH04E{'}Lj}L2RCMoH
RRRRRRRRRRRRFRRMEC_F_0#OOEC	RC8<F=RMEC_F_0#OOEC	RC8|CR0#C0_G;bs
RRRRRRRRRRRR8CM
RRRRRRRRCRRMR8
RRRRRCRRMR8
RRRRRCRRDR#CLHCoMH
`VV8CRpme_QQha _)tR
RRRRRRFRRMEC_F_0#OOEC	RC8<{=RI0H8E'{4L}j};C
`MV8H
RRRRRRRR8CMRR
RRRRRC
M8
RRRRORRFsPC_#0C0G_CbNs_DxD_C#sF:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRsRfF5#C00C#_bCGs=R=RH{I8{0E4j'L}R}22R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbNs_DxD_C#sFRPOFC8sC"
2;
RRRRORRFsPC_DND_CFM_0EF#E_OCCO	8R:
RRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	RFfs#FC5MEC_F_0#OOEC	RC8={=RI0H8E'{4L}4}2R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"DND_CFM_0EF#E_OCCO	8FROPCCs8;"2
RRRRMRC8/R/OMFsCOsRFsPCN
oCRRRRC
M8
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m




