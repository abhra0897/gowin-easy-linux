`ifndef ATCGPIO100_CONFIG_VH
`define ATCGPIO100_CONFIG_VH
`include "ae250_config.vh"
`include "ae250_const.vh"

//-------------------------------------------------
// GPIO Channel Number
//-------------------------------------------------
// Available value: 1~32
//`define ATCGPIO100_GPIO_NUM 32

//-------------------------------------------------
// GPIO Pull Option
//-------------------------------------------------
//`define ATCGPIO100_PULL_SUPPORT

//-------------------------------------------------
// GPIO Interrupt Option
//-------------------------------------------------
//`define ATCGPIO100_INTR_SUPPORT

//-------------------------------------------------
// GPIO Debounce Option
//-------------------------------------------------
//`define ATCGPIO100_DEBOUNCE_SUPPORT

`endif // ATCGPIO100_CONFIG_VH

