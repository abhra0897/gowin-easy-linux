@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)am_h B7mp"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
`RRHCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0MRC
RM`C8
HV
V`H8RCVm_ep1)]q B7_m
7 
IRRHRsCHOMN0CHP_DPN=M5HNHO0P=C=`pme_pqp_ mh142?':L44j'L;`

CHM8V/R/Rpme_q1])_ 7B m7
H
`VV8CRpme_1q1 _)am
h
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRFbsb0Cs$1Rq1a )_ mh_pBm7Z_X_
u;RRRR@b@5F8#CoOCRD
	2RRRR8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RRRR5f!5HM#k	IMFMC50#C0_G2bs2
2;RRRRCbM8sCFbs
0$RCR`MV8HRR//m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/eRmpB_X]i B_wmw
R
RbbsFC$s0R1q1 _)am_h B7mp_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R!fkH#MF	MI0M5C_#0CsGb2|2R-5>RRF5fMFCE005~C_#0CsGb2|2R|R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RR5NHMOP0HCRR<`pme_ mh_pBm7&2R&R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5#0C0G_Cb=sR=IR{HE80{NHMOP0HCN_PD2}}2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
2;RMRC8Fbsb0Cs$R

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)am_h B7mp_Ru:RNRR#s#C0sRbFsbC05$Rq 11)ma_hB _m_p7uR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFRMOF0MNH#FRlsFCRsCRD#0#RERNM4CR8NC##s80CR0LH#;"2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRqRR_1q1 _)am_h B7mp__XZuN:R#s#C0sRbFsbC05$Rq 11)ma_hB _m_p7XuZ_2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/Rpme_uQvpQQBaB_X]i B_wmw
M`C8RHV/m/ReXp_BB] iw_mwR

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRv1_q1a )_ mh_pBm7:_uRRRRNk##lbCRsCFbsR0$51q1 _)am_h B7mp_;u2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRvRR_1q1 _)am_h B7mp__XZuN:R#l#kCsRbFsbC05$Rq 11)ma_hB _m_p7XuZ_2R;
RM`C8RHV/m/ReQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/Rpme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_hR

RsRRCRoRr8IH04E-:Rj9F_MCO8FD#E_OCCO	8R;
RIRRHRsCr8IH04E-:Rj900C#_bCGsR_H=0R~C_#0CsGb;R
RRHRIsrCRI0H8E:-4j09RC_#0CsGb_4H_R0=RC_#0CsGb_-HRRI{{HE80-44{'}Lj}',4L;4}
C
oMNCs0
C
RRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRRHV5pme_eBm 1)_qahQYh_m2CRLoRHM:PRFDF_OP_Cs#HNM0
$
RRRROCFPsC_0#C0_G_bsOMENo
C:RRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25m5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRR!RRfN#0L5DC00C#_bCGs22R2R
RRRRRRRRRRRRRRRRRRDFP_POFC0s_5C"0#C0_G_bsOMENoOCRFsPCC28";R
RR8CMR#//N0MH$FROPNCso
C
RHRRVmR5eBp_m)e _)Bmh_ )mRh2LHCoMRR:F_PDOCFPsF_OssMC
R
RRDRNI#N$R5@@bCF#8RoCO2D	RoLCHRM
RRRRH5VR`pme_1)  1a_Qqthp=R!RL4'jL2RCMoH
RRRRHRRV5R500C#_bCGsRR^00C#_bCGs=2={8IH04E{'}Lj}L2RCMoH
RRRRRRRH5VR5NHMOP0HCm>`eqp_pmp_h2 1RR||5#0C0G_Cb=s!{8IH0HE{M0NOH_PCP}ND}R22LHCoMR
RRRRRRVRHR55!5#0C0G_CbHs_RR=={8IH04E{'}Lj}|2R|R
RRRRRRRRRRC50#C0_G_bsHRR&00C#_bCGs__H4!2R=IR{HE80{L4'j2}}2CRLo
HMRRRRRRRRRFRRMOC_F#D8_COEO8	CRR<=F_MCO8FD#E_OCCO	8RR|5C~0#C0_G2bs;R
RRRRRRMRC8R
RRRRRR8CM
RRRRCRRMR8
RRRRC
M8RRRRR#CDCCRLo
HM`8HVCmVReQp_h_Qa)
 tRRRRRMRFCF_OD_8#OOEC	RC8<{=RI0H8E'{4L}j};C
`MV8H
RRRRMRC8RR
RCRRM/8R/DRNI#N$
R
RRFROP_CsN_DDF_MCO8FD#E_OCCO	8R:
RORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	f2RsCF#5CFM_DOF8O#_E	COC=8R=IR{HE80{L4'42}}2R
RRRRRRRRRRRRRRRRRF_PDOCFPs5_0"DND_CFM_DOF8O#_E	COCO8RFsPCC28";R

RVRHRM5HNHO0P=CR=mR`eqp_pZp_ 1)m2CRLoRHM:PRFDF_OP_Cs00C#_bCGsD_NDC_xs
F#R
RRRRRROCFPsC_0#C0_G_bsN_DDxFCs#R:
RORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRfRRsCF#5#0C0G_Cb=sR=IR{HE80{NHMOP0HCN_PD2}}R
22RRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsD_NDC_xsRF#OCFPs"C82R;
RMRC8R

RVRHRM5HNHO0P=CR=mR`eqp_pmp_h2 1RoLCH:MRRDFP_POFC0s_C_#0CsGb_DND_CFM#R
R
RRRRPOFC0s_C_#0CsGb_DND_CFM#R:
RORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52RRm5`e)p_ a1 _t1QhRqp!4=R'2LjR
&&RRRRRRRRRRRRRRRRRfRRsCF#5#0C0G_Cb=sR=IR{HE80{NHMOP0HCN_PD2}}R
22RRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsD_NDM_FCO#RFsPCC28";R
RR8CM
CRRM/8R/sOFMRCsOCFPsCNo
MRC8C

MC8oMNCs0
C
`8CMH/VR/eRmpm_Be_ )m
h

