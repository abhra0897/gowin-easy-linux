`define DEF_AO_0_EN   
//`define DEF_AO_1_EN
//`define DEF_AO_2_EN
//`define DEF_AO_3_EN
//`define DEF_AO_4_EN
//`define DEF_AO_5_EN
//`define DEF_AO_6_EN
//`define DEF_AO_7_EN
//`define DEF_AO_8_EN
//`define DEF_AO_9_EN
//`define DEF_AO_10_EN
//`define DEF_AO_11_EN
//`define DEF_AO_12_EN
//`define DEF_AO_13_EN
//`define DEF_AO_14_EN
//`define DEF_AO_15_EN

// If CPU_0 sub-module is supported uncomment the following line
`define DBG_SUPPORTED_AO_0

// If CPU_1 sub-module is supported uncomment the following line
//`define DBG_SUPPORTED_AO_1

