@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ma_7u7_qa)QY
";
`RRHDMOkR8C"8#0_DFP_#0N	"3E
`

HCV8VeRmph_QQva_1Rt
RHRRMHH0NRD
RRRRRDFP_HHM0#_lo;_0RR//BDNDRC0ERCz#sCR7VCHM8MRQHv0RCN##o)CRFHk0M`C
CHM8V/R/m_epQahQ_tv1
H
`VV8CRpme_1q1 _)am
h
RsRbFsbC0q$R1)1 a7_m7q_u)YQa_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R^R55#0C0G_Cb2s2;R
RCbM8sCFbs
0$
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_7m7_)uqQ_aYXmZ_h _a1 a_X_u)uR;
RR@@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R5R5!H5f#	kMMMFI5#0C0G_Cb2s22
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRR_Rqq 11)ma_7u7_qa)QY:_uR#N#CRs0bbsFC$s0R15q1a )_7m7_)uqQ_aYuR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFM8#FCR0MFRECGH0LHR8F8RsbNH"0$2
;
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 a7_m7q_u)YQa__XZmah_ _1a )Xu_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)am_77uQq)aXY_Zh_m_1a aX_ uu)_2R
RRRRRRDRC#FCRPCD_sssF_"0500C#_bCGsFROMH0NMX#RRRFsZ;"2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRM
8
RRRRRmR`eqp_1v1z RR:LHCoMRR:F_PDNk##lRC
RRRRRvRR_1q1 _)am_77uQq)auY_:#RN#CklRFbsb0Cs$qR51)1 a7_m7q_u)YQa_;u2
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRvRR_1q1 _)am_77uQq)aXY_Zh_m_1a aX_ uu)_:R
RRRRRR#RN#CklRFbsb0Cs$qR51)1 a7_m7q_u)YQa__XZmah_ _1a )Xu_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_ho

CsMCN
0C
RRRRRHV5POFCosNCC_DPRCD!`=Rm_epB me)m_hhR 2LHCoMRR:F_PDOCFPsR
RRHRRVmR5eBp_m)e _h1qQ_aYmRh2LHCoMRR:F_PDOCFPsN_#M$H0
R
RRRRROCFPsC_0#C0_G_bsOMENo
C:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR!RRfN#0L5DC00C#_bCGs22RRR2
RRRRRRRRRRRRRRRRRFRRPOD_FsPC_"0500C#_bCGsE_ONCMoRPOFC8sC"
2;RRRRR8CMR#//N0MH$FROPNCsoRC
RCRRM
8
CoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
