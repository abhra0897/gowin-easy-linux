@ELDHs$NsR Q  S;SS
S
kR#CQ   371a_tpmQ4B_43ncN;DD
#
kC RQ 1 3ap7_mBtQ_Qq)aq]3pRp;RRRRRRRRR
R
kR#CQ   371a_tpmQzB_ht1Qh3 7q;pp
R
RRRRRRRRRRRRRRRRRRRRRRRRRR
R
b	NONRoCBumvmhh aH1R#R

R0RN0LsHkR0C#_$MLODN	F_LGL:RFCFDN;MR
R
RR0N0skHL0#CR$LM_D	NO_GLFRRFVBbFlFMMC0:#RRObN	CNoRRH#0Csk;R

R0RN0LsHkR0CLODN	F_LGN_b8H_bM#:R0MsHo
;
RNRR0H0sLCk0RM#$_bMFsCkMRL:RFCFDN
M;
RRRNs00H0LkCORG_blN:0R#soHM;R

R0RN0LsHkR0CGlO_NFbRVFRBlMbFC#M0Rb:RNNO	oHCR#DR"k;0"R-

-------------------------Xvz.----------------------------
--
B

mmvuha hRXvz.
R
RRRRuam)R
5
SRRRRRQj:MRHR8#0_oDFH
O;
RSRR4RQRH:RM0R#8F_Do;HO
R
SR1RRjRR:H#MR0D8_FOoH;S

RRRRmRR:FRk0#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFvVRzRX.:FRBlMbFCRM0H0#Rs;kC




-
-------------------------v.zX_apz6----------------------------
--
B

mmvuha hRXvz.z_pa
6R
RRRR)uma
R5
RSRRjRQRH:RM0R#8F_Do;HO
R
SRQRR4RR:H#MR0D8_FOoH;S

RRRR1:jRRRHM#_08DHFoO
;
SRRRR:mRR0FkR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apz6RR:BbFlFMMC0#RHRk0sC
;




-------------------------z-vXp._z-an-----------------------------



vBmu mhhvaRz_X.pnzaRR

RuRRmR)a5S

RRRRQ:jRRRHM#_08DHFoO
;
SRRRRRQ4:MRHR8#0_oDFH
O;
RSRRjR1RH:RM0R#8F_Do;HO
R
SRmRRRF:Rk#0R0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRan:FRBlMbFCRM0H0#Rs;kC




-
-------------------------v.zX_apz(----------------------------
--
B

mmvuha hRXvz.z_pa
(R
RRRR)uma
R5
RSRRjRQRH:RM0R#8F_Do;HO
R
SRQRR4RR:H#MR0D8_FOoH;S

RRRR1:jRRRHM#_08DHFoO
;
SRRRR:mRR0FkR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_apz(RR:BbFlFMMC0#RHRk0sC
;




-------------------------z-vXp._z-aU-----------------------------



vBmu mhhvaRz_X.pUzaRR

RuRRmR)a5S

RRRRQ:jRRRHM#_08DHFoO
;
SRRRRRQ4:MRHR8#0_oDFH
O;
RSRRjR1RH:RM0R#8F_Do;HO
R
SRmRRRF:Rk#0R0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvXp._zRaU:FRBlMbFCRM0H0#Rs;kC




-
-------------------------v.zX_XvzU----------------------------
--
B

mmvuha hRXvz.z_vX
UR
RRRR)uma
R5
RSRRjRQRH:RM0R#8F_Do;HO
R
SRQRR4RR:H#MR0D8_FOoH;S

RRRR1:jRRRHM#_08DHFoO
;
SRRRR:mRR0FkR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_XvzURR:BbFlFMMC0#RHRk0sC
;




-------------------------z-vXv._znX4-----------------------------
-

m
Bvhum Rhav.zX_Xvz4
nR
RRRR)uma
R5
RSRRjRQRH:RM0R#8F_Do;HO
R
SRQRR4RR:H#MR0D8_FOoH;S

RRRR1:jRRRHM#_08DHFoO
;
SRRRR:mRR0FkR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVv.zX_Xvz4:nRRlBFbCFMMH0R#sR0k
C;




------------------------v--z_X.vdzX.----------------------------
--
B

mmvuha hRXvz.z_vXRd.
R
RRmRu)5aR
R
SRQRRjRR:H#MR0D8_FOoH;S

RRRRQ:4RRRHM#_08DHFoO
;
SRRRRR1j:MRHR8#0_oDFH
O;
RSRRRRm:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvz.z_vXRd.:FRBlMbFCRM0H0#Rs;kC




-
-------------------------vczX-----------------------------
-

m
Bvhum RhavczXRR

RuRRmR)a5S

RRQj:MRHR8#0_oDFH
O;
QSR4RR:H#MR0D8_FOoH;S

RRQ.:MRHR8#0_oDFHRO;
R
SQ:dRRRHM#_08DHFoO
;
SjR1RH:RM0R#8F_Do;HO
R
S1:4RRRHM#_08DHFoO
;
SRRm:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzcRR:BbFlFMMC0#RHRk0sC
;




-------------------------z-vX-U-----------------------------



Bumvmhh azRvX
UR
RRRR)uma
R5
QSRjRR:H#MR0D8_FOoH;S

RRQ4:MRHR8#0_oDFH
O;
QSR.RR:H#MR0D8_FOoH;
R
SdRQRH:RM0R#8F_Do;HO
R
SQ:cRRRHM#_08DHFoO
;
S6RQRH:RM0R#8F_Do;HO
R
SQ:nRRRHM#_08DHFoO
;
S(RQRH:RM0R#8F_Do;HO
R
S1:jRRRHM#_08DHFoO
;
S4R1RH:RM0R#8F_Do;HO
R
S1:.RRRHM#_08DHFoO
;
SRRm:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzURR:BbFlFMMC0#RHRk0sC
;




-------------------------z-vX-4n----------------------------



Bumvmhh azRvXR4nRR

RuRRmR)a5S

RRQj:MRHR8#0_oDFH
O;
QSR4RR:H#MR0D8_FOoH;S

RRQ.:MRHR8#0_oDFHRO;
R
SQ:dRRRHM#_08DHFoO
;
ScRQRH:RM0R#8F_Do;HO
R
SQ:6RRRHM#_08DHFoO
;
SnRQRH:RM0R#8F_Do;HO
R
SQ:(RRRHM#_08DHFoO
;
SURQRH:RM0R#8F_Do;HO
R
SQ:gRRRHM#_08DHFoO
;
S4RQjRR:H#MR0D8_FOoH;S

R4Q4RH:RM0R#8F_Do;HO
R
SQR4.:MRHR8#0_oDFH
O;
QSR4:dRRRHM#_08DHFoO
;
S4RQcRR:H#MR0D8_FOoH;S

R6Q4RH:RM0R#8F_Do;HO
R
S1:jRRRHM#_08DHFoO
;
S4R1RH:RM0R#8F_Do;HO
R
S1:.RRRHM#_08DHFoO
;
SdR1RH:RM0R#8F_Do;HO
R
SmRR:FRk0#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFvVRznX4RB:RFFlbM0CMRRH#0Csk;



-

-------------------------Xvzd-.--------------------------
--
B

mmvuha hRXvzdR.R
R
RRmRu)5aR
R
SQ:jRRRHM#_08DHFoO
;
S4RQRH:RM0R#8F_Do;HO
R
SQ:.RRRHM#_08DHFoO
;R
QSRdRR:H#MR0D8_FOoH;S

RRQc:MRHR8#0_oDFH
O;
QSR6RR:H#MR0D8_FOoH;S

RRQn:MRHR8#0_oDFH
O;
QSR(RR:H#MR0D8_FOoH;S

RRQU:MRHR8#0_oDFH
O;
QSRgRR:H#MR0D8_FOoH;S

RjQ4RH:RM0R#8F_Do;HO
R
SQR44:MRHR8#0_oDFH
O;
QSR4:.RRRHM#_08DHFoO
;
S4RQdRR:H#MR0D8_FOoH;S

RcQ4RH:RM0R#8F_Do;HO
R
SQR46:MRHR8#0_oDFH
O;
QSR4:nRRRHM#_08DHFoO
;
S4RQ(RR:H#MR0D8_FOoH;S

RUQ4RH:RM0R#8F_Do;HO
R
SQR4g:MRHR8#0_oDFH
O;
QSR.:jRRRHM#_08DHFoO
;
S.RQ4RR:H#MR0D8_FOoH;S

R.Q.RH:RM0R#8F_Do;HO
R
SQ:.dRMRHR8#0_oDFH
O;
QSR.:cRRRHM#_08DHFoO
;
S.RQ6RR:H#MR0D8_FOoH;S

RnQ.RH:RM0R#8F_Do;HO
R
SQR.(:MRHR8#0_oDFH
O;
QSR.:URRRHM#_08DHFoO
;
S.RQgRR:H#MR0D8_FOoH;S

RjQdRH:RM0R#8F_Do;HO
R
SQRd4:MRHR8#0_oDFHRO;
R
S1:jRRRHM#_08DHFoO
;
S4R1RH:RM0R#8F_Do;HO
R
S1:.RRRHM#_08DHFoO
;
SdR1RH:RM0R#8F_Do;HO
R
S1:cRRRHM#_08DHFoO
;
SRRm:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRXvzd:.RRlBFbCFMMH0R#sR0k
C;




------------------------p--z-a4-----------------------------B

mmvuha hRapz4
R
RRRRt  h)RQB5hRQQ:aRR0LH_OPC0RFs:X=R"Rj"2
;
RRRRuam)R
5
SRRRR:wRR0FkR8#0_oDFH
O;
RRRRRRRRRQj:MRHR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;

0
N0LsHkR0C#_$MLODN	F_LGVRFRapz4RR:BbFlFMMC0#RHRk0sC
;
Ns00H0LkCORG_blNRRFVp4zaRO:RFFlbM0CMRRH#"0Dk"
;
S



-

-------------------------apz.----------------------------
-
Bumvmhh azRpa
.R
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=X""jR
2;
RRRR)uma
R5
RRRSRRRR:wRR0FkR8#0_oDFH
O;
RRRSRRRRRQj:MRHR8#0_oDFH
O;
RRRSRRRRRQ4:MRHR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;

N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:.RRlBFbCFMMH0R#sR0k
C;
0SN0LsHkR0CGlO_NFbRVzRpa:.RRlOFbCFMMH0R#DR"k;0"




-
-------------------------pdza-----------------------------
-
Bumvmhh azRpa
dR
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"j";R2
R
RRmRu)5aR
R
RRRSRRRRw:kRF00R#8F_Do;HO
R
RRRSRRjRQRH:RM0R#8F_Do;HO
R
RRRSRR4RQRH:RM0R#8F_Do;HO
R
RRRSRR.RQRH:RM0R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRapzdRR:BbFlFMMC0#RHRk0sC
;
S0N0skHL0GCRON_lbVRFRapzdRR:ObFlFMMC0#RHRk"D0
";




------------------------p--z-ac----------------------------
m
Bvhum RhapczaRR

RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjj";R2
R
RRmRu)5aR
R
RRRSRRRRw:kRF00R#8F_Do;HO
R
RRRSRRjRQRH:RM0R#8F_Do;HO
R
RRRSRR4RQRH:RM0R#8F_Do;HO
R
RRRSRR.RQRH:RM0R#8F_Do;HO
R
RRRSRRdRQRH:RM0R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRapzcRR:BbFlFMMC0#RHRk0sC
;
S0N0skHL0GCRON_lbVRFRapzcRR:ObFlFMMC0#RHRk"D0
";




------------------------p--z-a6----------------------------
m
Bvhum Rhap6zaRR

RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjj";R2
R
RRmRu)5aR
R
RRRSRRRRw:kRF00R#8F_Do;HO
R
RRRSRRjRQRH:RM0R#8F_Do;HO
R
RRRSRR4RQRH:RM0R#8F_Do;HO
R
RRRSRR.RQRH:RM0R#8F_Do;HO
R
RRRSRRdRQRH:RM0R#8F_Do;HO
R
RRRSRRcRQRH:RM0R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRapz6RR:BbFlFMMC0#RHRk0sC
;
S0N0skHL0GCRON_lbVRFRapz6RR:ObFlFMMC0#RHRk"D0
";




------------------------p--z-an----------------------------



Bumvmhh azRpa
nR
RRRRht  B)QRQ5RhRQa:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjRj"2
;
RRRRuam)R
5
RSRRRRRRwRR:FRk0#_08DHFoO
;
RSRRRRRRQ:jRRRHM#_08DHFoO
;
RSRRRRRRQ:4RRRHM#_08DHFoO
;
RSRRRRRRQ:.RRRHM#_08DHFoO
;
RSRRRRRRQ:dRRRHM#_08DHFoO
;
RSRRRRRRQ:cRRRHM#_08DHFoO
;
RSRRRRRRQ:6RRRHM#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFpVRzRan:FRBlMbFCRM0H0#Rs;kC
N
S0H0sLCk0R_GOlRNbFpVRzRan:FROlMbFCRM0H"#RD"k0;



-

-------------------------apz(----------------------------
-

m
Bvhum Rhap(zaRR

RtRR )h Q5BRRQQhaRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj";R2
R
RRmRu)5aR
R
RRRSRRRRw:kRF00R#8F_Do;HO
R
RRRSRRjRQRH:RM0R#8F_Do;HO
R
RRRSRR4RQRH:RM0R#8F_Do;HO
R
RRRSRR.RQRH:RM0R#8F_Do;HO
R
RRRSRRdRQRH:RM0R#8F_Do;HO
R
RRRSRRcRQRH:RM0R#8F_Do;HO
R
RRQRS6RR:H#MR0D8_FOoH;R

RRRSRQRRnRR:H#MR0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRpa:(RRlBFbCFMMH0R#sR0k
C;
0SN0LsHkR0CGlO_NFbRVzRpa:(RRlOFbCFMMH0R#DR"k;0"




-
-------------------------pUza-----------------------------



vBmu mhhpaRzRaU
R
RR RthQ )BRR5QahQRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR
2;
RRRR)uma
R5
RRRSRRRR:wRR0FkR8#0_oDFH
O;
RRRSRRRRRQj:MRHR8#0_oDFH
O;
RRRSRRRRRQ4:MRHR8#0_oDFH
O;
RRRSRRRRRQ.:MRHR8#0_oDFH
O;
RRRSRRRRRQd:MRHR8#0_oDFH
O;
RRRSRRRRRQc:MRHR8#0_oDFH
O;
RRRSRRRRRQ6:MRHR8#0_oDFH
O;
RRRSRRRRRQn:MRHR8#0_oDFH
O;
RRRSRRRRRQ(:MRHR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVpUzaRB:RFFlbM0CMRRH#0Csk;S

Ns00H0LkCORG_blNRRFVpUzaRO:RFFlbM0CMRRH#"0Dk"
;




-------------------------p-qz-------------------------------



Bumvmhh apRqz
R
RRRRt  h)RQB5
RR
RRRRRRRR7Rq7RR:Q hatR ):j=RR
;
RRRRRSRRRA1zRQ:Rhta  :)R=RR4;R

RRRRRRRRq177z:ARRaQh )t RR:=.
R;
RRRRRRRS RhRQ:Rhta  :)R=RRd;R

RRRRRRRSt: RRaQh )t RR:=c
R;
RSRRpRR RR:Q hatR ):6=R;R

RRRRRRRSBRzu:hRQa  t)=R:R;nR
R
RRRRRRBRR7:hRRaQh )t RR:=(
R;
RRRRRRRRzRBuhB7RQ:Rhta  :)R=;RU
R
SRRRRvazpRQ:Rhta  :)R=;Rg
R
SRRRRq_pzv m7RQ:Rhta  :)R=
Rj
RRRRS2;
R
RRmRu)5aR
R
S1Rzv:zRma0R#8F_Do;HO
R
SBamzRm:Rz#aR0D8_FOoH;
S
SjRQRQ:Rh0R#8F_Do;HO
R
SQR4:Q#hR0D8_FOoH;S

R:QdRRQh#_08DHFoO
;
SQRBhQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRqzRR:BbFlFMMC0#RHRk0sC
;




----------------------------7-ww-----------------------------



vBmu mhh7aRw
wR
RRRRht  B)QRQ5RhRQa:HRL0=R:R''j2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wRB:RFFlbM0CMRRH#0Csk;



-

-------------------------w-7w- ------------------------------
--
B

mmvuha hRw7w 
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
BSR RR:Q#hR0D8_FOoH;
S
SpRBiRR:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRwRw :FRBlMbFCRM0H0#Rs;kC




-
----------------------7--w-w1--------------------------------



Bumvmhh awR7w
1R
RRRRht  B)QRQ5Rh:QaR0LHRR:='R4'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
1SR :aRRRQh#_08DHFoO
;S
BSRp:iRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV71wwRB:RFFlbM0CMRRH#0Csk;



-

-------------------------7--w w1-------------------------------------
-

m
Bvhum Rha71ww 
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
1SR :aRRRQh#_08DHFoO
;
S RB:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7w1: RRlBFbCFMMH0R#sR0k
C;




------------------------w7w)--------------------------------
--
B

mmvuha hRw7w)
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
)SR a1 RQ:Rh0R#8F_Do;HOSS

RiBpRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:)RRlBFbCFMMH0R#sR0k
C;




---------------------------7)ww ------------------------------------
-

m
Bvhum Rha7)ww 
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
)SR a1 RQ:Rh0R#8F_Do;HO
R
SBR :Q#hR0D8_FOoH;
S
SpRBiRR:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRw w)RB:RFFlbM0CMRRH#0Csk;



-

-------------------------7--w-wu-------------------------------------
-

m
Bvhum Rha7uwwRR

RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
S)Ru a1 :hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wuRR:BbFlFMMC0#RHRk0sC
;




-------------------------w-7w-u --------------------------------------------



Bumvmhh awR7wRu 
R
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R u)1R a:hRQR8#0_oDFH
O;
BSR Q:Rh0R#8F_Do;HOSS

RiBpRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRu :FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--w-wB-----------------------------
--
B

mmvuha hRw7wB
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
BSRp) qRQ:Rh0R#8F_Do;HOSS

RiBpRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w:BRRlBFbCFMMH0R#sR0k
C;




----------------------------w-7w-B -----------------------------------------
-

m
Bvhum Rha7Bww 
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
BSRp) qRQ:Rh0R#8F_Do;HO
R
SBR :Q#hR0D8_FOoH;
S
SpRBiRR:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRw wBRB:RFFlbM0CMRRH#0Csk;



-

-------------------------w7wh----------------------------
--
B

mmvuha hRw7wh
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='2j';
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;S
BSRp:iRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7hwwRB:RFFlbM0CMRRH#0Csk;



-

-----------------w7wh- ------------------------------
--
B

mmvuha hRw7wh
 R
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
R
RRmRu)5aR
R
STRR:mRza#_08DHFoO
;S
7SRRQ:Rh0R#8F_Do;HO
R
SB: RRRQh#_08DHFoO
;S
BSRp:iRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww RR:BbFlFMMC0#RHRk0sC
;




-------------------------w7wh-1------------------------------
--
B

mmvuha hRw7wh
1R
RRRRht  B)QRQ5Rh:QaR0LHRR:='R4'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
1SR :aRRRQh#_08DHFoO
;S
BSRp:iRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww1RR:BbFlFMMC0#RHRk0sC
;




----------------------------7hww1- -------------------------------------



Bumvmhh awR7w h1RR

RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
S R1aRR:Q#hR0D8_FOoH;S

R:B RRQh#_08DHFoO
;S
BSRp:iRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7hww1: RRlBFbCFMMH0R#sR0k
C;




----------------------------w-7w-h)---------------------------------



vBmu mhh7aRw)whRR

RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
S R)1R a:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:)RRlBFbCFMMH0R#sR0k
C;




---------------------------7hww)- ----------------------------------
--
B

mmvuha hRw7whR) 
R
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R1)  :aRRRQh#_08DHFoO
;
S RB:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whR) :FRBlMbFCRM0H0#Rs;kC




-
--------------------------w-7w-hu-------------------------------------
-

m
Bvhum Rha7hwwu
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='R4'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
uSR)  1aQ:Rh0R#8F_Do;HOSS

RiBpRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7wRhu:FRBlMbFCRM0H0#Rs;kC




-
-------------------------7hwwu- ------------------------------------------
--
B

mmvuha hRw7whRu 
R
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R u)1R a:hRQR8#0_oDFH
O;
BSR Q:Rh0R#8F_Do;HOSS

RiBpRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVwR7w huRB:RFFlbM0CMRRH#0Csk;



-

----------------------------7hwwB--------------------------------------------



vBmu mhh7aRwBwhRR

RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
SpRB Rq):hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7wh:BRRlBFbCFMMH0R#sR0k
C;




----------------------------w-7w hB-----------------------------------------
--
B

mmvuha hRw7whRB 
R
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R Bpq:)RRRQh#_08DHFoO
;
S RB:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRw7whRB :FRBlMbFCRM0H0#Rs;kC




-
------------------------------p-7-----------------------------------------
-

m
Bvhum Rha7
pR
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
R
RRmRu)5aR
R
STRR:mRza#_08DHFoO
;S
7SRRQ:Rh0R#8F_Do;HOSS

R:tRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7:pRRlBFbCFMMH0R#sR0k
C;




------------------------p-7 -----------------------------------



Bumvmhh apR7 
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
BSR Q:Rh0R#8F_Do;HOSS

R:tRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rp :FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--p-B----------------------------------
-

m
Bvhum Rha7RpB
R
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R Bpq:)RRRQh#_08DHFoO
;S
tSRRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVpR7BRR:BbFlFMMC0#RHRk0sC
;




-----------------------------B7p ------------------------------------



vBmu mhh7aRpRB 
R
RR RthQ )BRR5QahQRL:RH:0R=jR'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R Bpq:)RRRQh#_08DHFoO
;S
tSRRQ:Rh0R#8F_Do;HO
R
SBR :Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRB :FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--p-u----------------------------------
-

m
Bvhum Rha7Rpu
R
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:#_08DHFoO
;
S)Ru a1 RQ:Rh0R#8F_Do;HOSS

RRt:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:uRRlBFbCFMMH0R#sR0k
C;




----------------------------p-7u- ----------------------------------
-

m
Bvhum Rha7 puRR

RtRR )h Q5BRRQQhaRR:LRH0:'=R42'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
S)Ru a1 RQ:Rh0R#8F_Do;HOSS

R:tRRRQh#_08DHFoO
;
S RB:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRu7p RR:BbFlFMMC0#RHRk0sC
;




------------------------7-ph-----------------------------------------



vBmu mhh7aRp
hR
RRRRht  B)QRQ5RhRQa:HRL0=R:R''jRS2;
R
RRmRu)5aR
R
STRR:mRza#_08DHFoO
;S
7SRRQ:Rh0R#8F_Do;HOSS

R:tRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7Rph:FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--p-h ---------------------------------
-

m
Bvhum Rha7 phRR

RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
S RB:hRQR8#0_oDFHSO;
R
StRR:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRh :FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--p-hB---------------------------------
--
B

mmvuha hRh7pB
R
RRRRt  h)RQB5hRQQ:aRR0LHRR:='Rj'2
;S
RRRR)uma
R5
TSRRm:Rz#aR0D8_FOoH;
S
SRR7:hRQR8#0_oDFH
O;
BSRp) qRQ:Rh0R#8F_Do;HOSS

R:tRRRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7BphRB:RFFlbM0CMRRH#0Csk;



-

----------------------------7Bph ------------------------------------



vBmu mhh7aRp hBRR

RtRR )h Q5BRRQQhaRR:LRH0:'=Rj2'R;
S
RRRRuam)R
5
SRRT:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
SpRB Rq):hRQR8#0_oDFHSO;
R
StRR:Q#hR0D8_FOoH;S

R:B RRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7Bph RR:BbFlFMMC0#RHRk0sC
;




-----------------------------h7pu------------------------------------



vBmu mhh7aRpRhu
R
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:#_08DHFoO
;
S)Ru a1 RQ:Rh0R#8F_Do;HOSS

RRt:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRpRhu:FRBlMbFCRM0H0#Rs;kC




-
--------------------------7--p hu------------------------------------



Bumvmhh apR7hRu 
R
RR RthQ )BRR5QahQRL:RH:0R=4R'';R2SR

RuRRmR)a5S

R:TRRamzR8#0_oDFHSO;
R
S7RR:Q#hR0D8_FOoH;S

R u)1R a:hRQR8#0_oDFHSO;
R
StRR:Q#hR0D8_FOoH;S

R:B RRQh#_08DHFoOR

R2RR;
S
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7uph RR:BbFlFMMC0#RHRk0sC
;




-----------------eQh---------------------------------



vBmu mhhQaRh
eR
RRRR)uma
R5
RRRRmSRRm:Rz#aR0D8_FOoH;R

RSRRR:QRRRQh#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVRh:eRRlBFbCFMMH0R#sR0k
C;








--------------------Q--A-zw------------------------------------



Bumvmhh aARQz
wR
RRRR)uma
R5
RRRRmSRRm:Rz#aR0D8_FOoH;R

RSRRR:QRRRQh#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVRARzw:FRBlMbFCRM0H0#Rs;kC




-
-----------------------------mwAz-------------------------------------
--
B

mmvuha hRzmAw
R
RRRRuam)R
5
RRRRSRRm:zRma0R#8F_Do;HO
R
RRRRSQRR:Q#hR0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVARmz:wRRlBFbCFMMH0R#sR0k
C;




------------------------------------zaAw---------------------------



Bumvmhh aARaz
wR
RRRR)uma
R5
RRRRRSm:zRma0R#8F_Do;HO
R
RRQRSRQ:Rh0R#8F_Do;HO
R
RRmRS :hRRRQh#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFaVRARzw:FRBlMbFCRM0H0#Rs;kC
R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRzaAwRR:BbFlFMMC0#RHR""m;







----------------------------AQmz-w------------------------------
-

m
Bvhum RhaQzmAw
R
RRRRuam)R
5
RRRRSRmR:zRmaRRR#_08DHFoO
;
RRRRSRQm:hRQmRza#_08DHFoO
;
RRRRRRSQRQ:RhRRRR8#0_oDFH
O;
RSRR RmhRR:QRhRR0R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRAQmz:wRRlBFbCFMMH0R#sR0k
C;




--------------------------------7-Q7-)-------------------------



Bumvmhh a7RQ7
)R
RRRRht  B)QR
5
S_TjQahQRL:RH:0R=jR''
;
S_T4QahQRL:RH:0R=jR''R

R2RR;
S
RRRRuam)R
5
SjRTRm:Rz#aR0D8_FOoH;S

RRT4:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
SpRBiQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV7RQ7:)RRlBFbCFMMH0R#sR0k
C;




--------------------------------7-Q7-)B-------------------------
-

m
Bvhum RhaQ)77B
R
RRRRt  h)RQB5
R
S_TjQahQRL:RH:0R=jR''
;
S_T4QahQRL:RH:0R=jR''R

R2RR;
S
RRRRuam)R
5
SjRTRm:Rz#aR0D8_FOoH;S

RRT4:zRma0R#8F_Do;HOSS

R:7RRRQh#_08DHFoO
;
SpRB :q)RRQh#_08DHFoO
;S
BSRpRi:Q#hR0D8_FOoH
R
RR;R2SC

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVR7B7)RB:RFFlbM0CMRRH#0Csk;







-------------------------------m)77---------------------
-

m
Bvhum Rham)77RR

RtRR )h Q5BRRR

RRRRRaRRXiBp_pumRL:RH:0R=jR''-;-':j')HH#MCoR8RoCFbk0kR0;':4'wDNDHRMoCC8oR0FkbRk0RRRRR
RR
RRRRRRRRhBm1haqahRQQ:aRR8#0_oDFH:OR=jR''
R
RRRR2
;S
RRRR)umaRR5
R
SRTRRjRR:mRza#_08DHFoO
;S
RSRR4RTRm:Rz#aR0D8_FOoH;
S
SRRRRR7j:hRQR8#0_oDFH
O;
RSRR4R7RQ:Rh0R#8F_Do;HO
R
SRaRRXRR:Q#hR0D8_FOoH;S

RRRRBRpi:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR7m7)RR:BbFlFMMC0#RHRk0sC
;





-
------------------------------7m7)-B---------------------
m
Bvhum Rham)77B
R
RRRRt  h)RQB5
R
RRRRRRRRapXBim_upRR:LRH0:'=Rj-';-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bkRRRRRRRR
R
RRRRRRmRBhq1ahQaRhRQa:0R#8F_DoRHO:'=Rj
'R
RRRRS2;
R
RRmRu)5aR
R
ST:jRRamzR8#0_oDFHSO;
R
ST:4RRamzR8#0_oDFHSO;
R
S7:jRRRQh#_08DHFoO
;
S4R7RQ:Rh0R#8F_Do;HOSS

RRaX:hRQR8#0_oDFHSO;
R
SBRpi:hRQR8#0_oDFH
O;
BSRp) q:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR7m7):BRRlBFbCFMMH0R#sR0k
C;




-

----------------------------------------Q17 c-------------------------------



Bumvmhh a7RQ R1c
t
S )h Q5BR
S
St 1)hRR:#H0sM:oR=VR"NCD#"
;
S1Sp)R h:0R#soHMRR:="k0sC
"
S
2;
mSu)5aR
S
S7RR:Q#hR0D8_FOoH;S

SpBqQ:ARRRQh#_08DHFoO
;
S S)1R a:hRQR8#0_oDFH
O;
wSSBRpi:hRQR8#0_oDFH
O;
uSSBRpi:hRQR8#0_oDFH
O;
TSSjRR:mRza#_08DHFoO
;
S4STRm:Rz#aR0D8_FOoH;S

SRT.:zRma0R#8F_Do;HO
S
ST:dRRamzR8#0_oDFH
O
S
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR Q71:cRRlBFbCFMMH0R#sR0k
C;




-

---------------------------------Q--e Q7m-------------------------------



Bumvmhh aeRQQm7 RR

RtRR )h Q5BR
S
St 1)hRR:#H0sM:oR=VR"NCD#"
;
S1Sp)R h:0R#soHMRR:="k0sC
"
RRRR2
;
RRRRuam)R
5
SRS7:hRQR8#0_oDFH
O;
)SS a1 RQ:Rh0R#8F_Do;HO
S
SBQqpARR:Q#hR0D8_FOoH;S

SpwBiRR:Q#hR0D8_FOoH;S

SpuBiRR:Q#hR0D8_FOoH;S

SRTj:zRma0R#8F_Do;HO
S
ST:4RRamzR8#0_oDFH
O;
TSS.RR:mRza#_08DHFoO
;
SdSTRm:Rz#aR0D8_FOoH;S

SRTc:zRma0R#8F_Do;HO
S
ST:6RRamzR8#0_oDFH
O;
TSSnRR:mRza#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVRe Q7mRR:BbFlFMMC0#RHRk0sC
;




---------------------------------Q--7U 1-------------------------------------



vBmu mhhQaR7U 1RR

RtRR )h Q5BR
R
SRtRR1h) R#:R0MsHo=R:RN"VD"#C;S

S)p1 :hRRs#0HRMo:"=R0Csk"R

R2RR;R

RuRRmR)a5S

S)7, a1 RQ:Rh0R#8F_Do;HO
S
SBQqpARR:Q#hR0D8_FOoH;S

SpwBiB,up:iRRRQh#_08DHFoO
;
SjSTRm:Rz#aR0D8_FOoH;S

SRT4:zRma0R#8F_Do;HO
S
ST:.RRamzR8#0_oDFH
O;
TSSdRR:mRza#_08DHFoO
;
ScSTRm:Rz#aR0D8_FOoH;S

SRT6:zRma0R#8F_Do;HO
S
ST:nRRamzR8#0_oDFH
O;
TSS(RR:mRza#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVR7U 1RB:RFFlbM0CMRRH#0Csk;







------------------------------------Q--74 1j--------------------------------
--
B

mmvuha hR Q71R4j
R
RR RthQ )B
R5
RSRR1Rt)R h:0R#soHMRR:="DVN#;C"
S
Sp 1)hRR:#H0sM:oR=0R"s"kC
R
RR;R2
R
RRmRu)5aR
S
S7 ,)1R a:hRQR8#0_oDFH
O;
BSSqApQRQ:Rh0R#8F_Do;HO
S
SwiBp,puBiRR:Q#hR0D8_FOoH;S

SRTj:zRma0R#8F_Do;HO
S
ST:4RRamzR8#0_oDFH
O;
TSS.RR:mRza#_08DHFoO
;
SdSTRm:Rz#aR0D8_FOoH;S

SRTc:zRma0R#8F_Do;HO
S
ST:6RRamzR8#0_oDFH
O;
TSSnRR:mRza#_08DHFoO
;
S(STRm:Rz#aR0D8_FOoH;S

SRTU:zRma0R#8F_Do;HO
S
ST:gRRamzR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVQ17 4:jRRlBFbCFMMH0R#sR0k
C;




-

------------------------m)1 c----------------------------
--
B

mmvuha hR m1)
cR
 SthQ )B
R5
tSS1h) R#:R0MsHo=R:RN"VD"#C;S

S)p1 :hRRs#0HRMo:"=R0Csk"
;
RRRRRRRR]RWp:0R#soHMRR:="DVN#;C"-0-"s"kC;VR"NCD#"R

RRRRRaRRXiBp_pumRL:RH:0R=jR'''--j)':HM#Ho8RCoFCRkk0b0';R4w':NHDDMCoR8RoCFbk0k
0
S
2;
mSu)5aR
S
S7:jRRRHM#_08DHFoO
;
S4S7RH:RM0R#8F_Do;HO
S
S7:.RRRHM#_08DHFoO
;
SdS7RH:RM0R#8F_Do;HO
S
SaRXj:MRHR8#0_oDFH
O;
aSSX:4RRRHM#_08DHFoO
;
SBSup:iRRRHM#_08DHFoO
;
S S)1R a:MRHR8#0_oDFH
O;
wSSBRpi:MRHR8#0_oDFH
O;
TSSjRR:mRza#_08DHFoO
;
S4STRm:Rz#aR0D8_FOoH
2
S;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFmVR1c )RB:RFFlbM0CMRRH#0Csk;







--------------------Qme7- m---------------------------------



vBmu mhhmaRe Q7m
R
Sht  B)Q5S

S)t1 :hRRs#0HRMo:"=RV#NDC
";
pSS1h) R#:R0MsHo=R:Rs"0k
C"
;S2
u
SmR)a5S

SR7j:MRHR8#0_oDFH
O;
7SS4RR:H#MR0D8_FOoH;S

SR7.:MRHR8#0_oDFH
O;
7SSdRR:H#MR0D8_FOoH;S

SR7c:MRHR8#0_oDFH
O;
7SS6RR:H#MR0D8_FOoH;S

SR7n:MRHR8#0_oDFH
O;
uSSBRpi:MRHR8#0_oDFH
O;
)SS a1 RH:RM0R#8F_Do;HO
S
SwiBpRH:RM0R#8F_Do;HO
S
STRR:mRza#_08DHFoOS

2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVm7eQ :mRRlBFbCFMMH0R#sR0k
C;




-------------------- m1)-U----------------------------------



vBmu mhhmaR1U )RR

RtRR )h Q5BR
R
RRtRS1h) R#:R0MsHo=R:RN"VD"#C;R

RSRRp 1)hRR:#H0sM:oR=0R"s"kC;R

RRRRR]RRW:pRRs#0HRMo:"=RV#NDC
";
RRRRRRRRBaXpui_m:pRR0LHRR:='-j'-''j:#)HHRMoCC8oR0Fkb;k0R''4:DwNDoHMRoC8CkRF00bk
R
RR;R2
R
RRmRu)5aR
R
RRRRRRjS7RH:RM0R#8F_Do;HO
R
RRRRRR4S7RH:RM0R#8F_Do;HO
R
RRRRRR.S7RH:RM0R#8F_Do;HO
R
RRRRRRdS7RH:RM0R#8F_Do;HO
R
RRRRRRcS7RH:RM0R#8F_Do;HO
R
RRRRRSR76:MRHR8#0_oDFH
O;
RRRRRRRSR7n:MRHR8#0_oDFH
O;
RRRRRRRSR7(:MRHR8#0_oDFH
O;
RRRRRRRSjaXRH:RM0R#8F_Do;HO
R
RRaRSX:4RRRHM#_08DHFoO
;
SRRRR.aXRH:RM0R#8F_Do;HO
R
SRaRRX:dRRRHM#_08DHFoO
;
SRRRRpuBiRR:H#MR0D8_FOoH;S

RRRR)  1aRR:H#MR0D8_FOoH;S

RRRRwiBpRH:RM0R#8F_Do;HO
R
RRRRRRjSTRm:Rz#aR0D8_FOoH;R

RRRRRTRS4RR:mRza#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFmVR1U )RB:RFFlbM0CMRRH#0Csk;







-------------------- m1)-4j---------------------------------
-
Bumvmhh a1Rm j)4RS

t  h)RQB5S

S)t1 :hRRs#0HRMo:"=RV#NDC
";
pSS1h) R#:R0MsHo=R:Rs"0k
C"
;S2
u
SmR)a5S

SR7j:MRHR8#0_oDFH
O;
7SS4RR:H#MR0D8_FOoH;S

SR7.:MRHR8#0_oDFH
O;
7SSdRR:H#MR0D8_FOoH;S

SR7c:MRHR8#0_oDFH
O;
7SS6RR:H#MR0D8_FOoH;S

SR7n:MRHR8#0_oDFH
O;
7SS(RR:H#MR0D8_FOoH;S

SR7U:MRHR8#0_oDFH
O;
7SSgRR:H#MR0D8_FOoH;S

SpuBiRR:H#MR0D8_FOoH;S

S1)  :aRRRHM#_08DHFoO
;
SBSwp:iRRRHM#_08DHFoO
;
SRST:zRma0R#8F_Do
HO
;S2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rm j)4RB:RFFlbM0CMRRH#0Csk;







-

-----------------Q--mp7 q-Y----------------------------------



vBmu mhhQaRmp7 q
YR
 SthQ )BRR5R1B_aQqaBp_7YRR:HCM0oRCs:j=R2-;-R4j~.
(
S)uma
R5
7SSQRR:Q#hR0D8_FOoH;S

Sa17q:uRRRQh#_08DHFoO
;
S S1a:hRRRQh#_08DHFoO
;
SqSepRz :hRQR8#0_oDFH
O;
7SSmRR:mRza#_08DHFoO
;
SwS7Rm:Rz#aR0D8_FOoH
2
S;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFQVRmp7 q:YRRlBFbCFMMH0R#sR0k
C;




--------------------vQ ---------------------------------
-

m
Bvhum RhaQR v
t
S )h Q
B5
WSSQQh1Z: RRs#0HRMo:"=R1pvqp
";
tSS1h) R#:R0MsHo=R:RN"VD"#C;S

S)p1 :hRRs#0HRMo:"=R0Csk"S

2
;
S)uma
R5
7SSRH:RM0R#8F_Do;HO
S
SBRpi:MRHR8#0_oDFH
O;
)SS a1 RH:RM0R#8F_Do;HO
S
SviBp:MRHR8#0_oDFH
O;
pSSq:tRR0FkR8#0_oDFH
O;
pSS Rq7:kRF00R#8F_Do
HO
;S2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV RQvRR:BbFlFMMC0#RHRk0sC
;





-
-------------------1u-------------------------------------
-
Bumvmhh auR1RR

RtRR )h Q5BR
R
SA_QaWaQ7]RR:HCM0oRCs:.=d;R--4.,R,,RcRRU,4Rn,d
.
S R)qv7_mR7 :HRL0=R:R''j;R--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
R
SWa)Q m_v7: RR0LH_OPC0RFs:"=Rj;j"-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8
C
RRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"-Y-1hRB,qh1YBS

RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
R
RR;R2
R
RRmRu)5aR
R
S7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
R
SB,piR,B m,B )  1a),W RR:H#MR0D8_FOoH;S

RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;
RRRRASRp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
R
S7:QRRRHM#_08DHFoOC_POs0F5Rd48MFI0jFR2R

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF1VRuRR:BbFlFMMC0#RHRk0sC
;





-
--------------------------u-1X-g--------------------------------------B

mmvuha hRX1ug
R
RRRRt  h)RQB5
R
SQRAaQ_W7Ra]:MRH0CCos=R:g
;
S R)qv7_mR7 :HRL0=R:R''j;R--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
R
SWa)Q m_v7: RR0LH_OPC0RFs:j="j-";-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCS

RiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"-Y-1hRB,qh1YBS

RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
R
RR;R2
R
RRmRu)5aR
R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
R
SB,piR,B m,B )  1a),W RR:H#MR0D8_FOoH;S

RRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;
7SRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj;R

RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj



RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV1guXRB:RFFlbM0CMRRH#0Csk;







-

---------------------------------u17A---------------------------------------
m
Bvhum Rha1A7uRR

RtRR )h Q5BRRS

RRRRA_QaWaQ7]R_j:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.S

RRRRA_QaWaQ7]R_4:MRH0CCos=R:4Rn;-4-R,,R.RRc,U4,Rnd,R.S

RRRR)7 q_7vm RR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8C
RRRRRRRRiAp_p1 _:jRR0LH_OPC0RFs:"=Rj"jj;R

RRRRRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBS

RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
R
RR;R2
R
RRmRu)5aR
R
SR7RRmRR:FRk0#_08DHFoOC_POs0F5Rd48MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,.
2;
RSRRpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1a:ARRRHM#_08DHFoO
;
SRRRRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
R
RRRRRRpRAip1 qp,Aip1 ARR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
R
SR7RRQRR:H#MR0D8_FOoH_OPC05Fsd84RF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV7R1u:ARRlBFbCFMMH0R#sR0k
C;
-

---------------------------------u17X-gA-------------------------------------
-
Bumvmhh a7R1uAXgRR

RtRR )h Q5BRRS

RRRRA_QaWaQ7]R_j:MRH0CCos=R:4RU;-g-R,UR4,nRd
R
SRARRQWa_Q]7a_:4RR0HMCsoCR4:=U-;R-,RgR,4UR
dn
RSRR R)qv7_mR7 :HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCS

RRRRA_pi1_ pjRR:L_H0P0COF:sR=jR"j;j"
R
SRARRp1i_ 4p_RL:RHP0_CFO0s=R:Rj"jj
";
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YBR";-Y-1hRB,qh1YBS

RRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRR
R
RRRR2
;
RRRRuam)R
5
SRRRRR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;S

RRRRBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A aRH:RM0R#8F_Do;HO
R
SRqRR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2
;
RRRRRRRRA1pi ,pqA1pi RpA:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2
;
SRRRRR7Q:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV1X7ug:ARRlBFbCFMMH0R#sR0k
C;
-

-------------------------7--u-A--------------------------------------



vBmu mhh7aRu
AR
RRRRht  B)QR
5
SASRQWa_Q]7a_:jRR0HMCsoCR4:=n
;R
RSSA_QaWaQ7]R_4:MRH0CCos=R:4Rn;
S
SRq) 7m_v7R j:HRL0=R:R''j;-R-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCS

S R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
SWSR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"RR--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8C
RSSWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
R
RRRRSA_pi1_ pjRR:L_H0P0COF:sR=jR"j;j"
R
RRRRSA_pi1_ p4RR:L_H0P0COF:sR=jR"j;j"
R
RRRRRR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;-R-1BYh,1RqY
hB
RSSQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
"
RRRR2
;
RRRRuam)R
5
S7SRm7q,m:ARR0FkR8#0_oDFHPO_CFO0s654RI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5j4;n2
S
SRiBpqp,BiRA,B, qB, AmqB , mBA ,)1q a,1)  ,aAWq) , W)ARR:H#MR0D8_FOoH;S

S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R

RSRRRiAp1q p,iAp1A pRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;
RSS7,Qq7RQA:MRHR8#0_oDFHPO_CFO0s654RI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV7RuA:FRBlMbFCRM0H0#Rs;kC



----------------------------7guXA---------------------------------------
m
Bvhum Rha7guXA
R
RRRRt  h)RQB5
R
SRRRRaAQ_7WQaj]_RH:RMo0CC:sR=;4URR--g4,RUS

RRRRA_QaWaQ7]R_4:MRH0CCos=R:4RU;-g-R,UR4
R
SR)RR _q7v m7jRR:LRH0:'=RjR';-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8C
RSRR R)qv7_m47 RL:RH:0R=jR''-;R-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
SRRRRQW)av _mj7 RL:RHP0_CFO0s=R:Rj"j"-;R-jRj:FRMsDlNR8lFCj;R4I:RsCH0-s0EFEkoR8lFC4;Rjs:RC-N8LFCVsIC-sCH0R8lFCS

RRRRWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;-R-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
R
RRRRRRpRAi _1pR_j:HRL0C_POs0FRR:="jjj"
;
RRRRRRRRA_pi1_ p4RR:L_H0P0COF:sR=jR"j;j"
R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1h
B
SRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
R
RRRR2
;
RRRRuam)R
5
SRRRRq7m,A7mRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2RjRR:=OPFM_8#0_oDFHPO_CFO0s,5j4;U2
R
SRBRRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;
RSRR7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;S

RRRR7RQq:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;
RRRRRRRRiAp1q p,iAp1A pRH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;
RSRRQR7ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR7XRgA:FRBlMbFCRM0H0#Rs;kC








-
---------------------------------1-7u-------------------------------------
-

m
Bvhum Rha1R7u
R
RR RthQ )BRR5
R
SA_QaWaQ7]R_j:MRH0CCos=R:4-n;-,R4RR.,cU,R,nR4,.Rd
R
SA_QaWaQ7]R_4:MRH0CCos=R:4-n;-,R4RR.,cU,R,nR4,.Rd
R
S)7 q_7vm RR:LRH0:'=Rj-';-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
RRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";
RRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"-Y-1hRB,qh1YBS

RQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v4_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v6_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vg_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v7_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRR
R
RR;R2
R
RRmRu)5aR
R
S7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
R
SBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A a, W)q),W :ARRRHM#_08DHFoO
;
S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R

RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;S

RR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV1R7u:FRBlMbFCRM0H0#Rs;kC







---------------------------------7-1u-Xg-------------------------------------
-
Bumvmhh a7R1uRXg
R
RR RthQ )BRR5
R
SA_QaWaQ7]R_j:MRH0CCos=R:4-U;-,RgR,4UR
dn
ASRQWa_Q]7a_:4RR0HMCsoCR4:=U-;-RRg,4RU,d
n
S R)qv7_mR7 :HRL0=R:R''j;R--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
R
SA_pi1R p:HRL0C_POs0FRR:="jjj"
;
RRRRR1)  va_mR7 :0R#soHMRR:="h1YB-";-h1YBq,R1BYh
R
SQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rj :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4 :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R..:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.n:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.q:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R. :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd.:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdn:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdq:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rd :HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRRR

R2RR;R

RuRRmR)a5S

RR7m:kRF00R#8F_Do_HOP0COFds56FR8IFM0R:j2=MOFP0_#8F_Do_HOP0COFjs5,2dn;S

RiBpqp,BiRA,B, qB, Am,B )  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2
;
RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2
;
SQR7RH:RM0R#8F_Do_HOP0COFds56FR8IFM0R
j2
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRu17X:gRRlBFbCFMMH0R#sR0k
C;




-

-------------------------7--u---------------------------------------



Bumvmhh auR7RR

RtRR )h Q5BR
S
SRaAQ_7WQaj]_RH:RMo0CC:sR=;4nRS

SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;
R
S)SR _q7v m7jRR:LRH0:'=Rj-';-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
S)SR _q7v m74RR:LRH0:'=Rj-';-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
SWSR) Qa_7vm :jRR0LH_OPC0RFs:"=Rj;j"-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8
C
SWSR) Qa_7vm :4RR0LH_OPC0RFs:"=Rj;j"-j-RjM:RFNslDFRl8RC;jR4:I0sHCE-0soFkEFRl8RC;4Rj:s8CN-VLCF-sCI0sHCFRl8
C
RRRRSpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
R
RRRRRR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;1--Y,hBRYq1h
B
SQSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SQSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSSQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
S
SRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"R

R2RR;R

RuRRmR)a5S

SmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R468MFI0jFR2O:=F_MP#_08DHFoOC_POs0F54j,n
2;
RSSBqpi,iBpAB,R Bq, mA,B, qmAB ,1)  ,aq)  1aWA,), qWA) RH:RM0R#8F_Do;HO
S
SRqq7,Aq7RH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2
R
RRRRSA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;S

SQR7qQ,7ARR:H#MR0D8_FOoH_OPC05Fs486RF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVuR7RB:RFFlbM0CMRRH#0Csk;







----------------------------X7ug---------------------------------------
m
Bvhum Rha7guXRR

RtRR )h Q5BRRS

RaAQ_7WQaj]_RH:RMo0CC:sR=;4U-g-R,UR4
R
SA_QaWaQ7]R_4:MRH0CCos=R:4-U;-,RgR
4U
)SR _q7v m7jRR:LRH0:'=Rj-';-:RjRbL$NR##lCF8;:R4RbbHCMDHCFRl8
C
S R)qv7_m47 RL:RH:0R=jR''-;-RRj:LN$b#l#RF;8CRR4:bCHbDCHMR8lFCS

RQW)av _mj7 RL:RHP0_CFO0s=R:Rj"j"-;-R:jjRsMFlRNDlCF8;4Rj:sRIH-0C0FEskRoElCF8;jR4:CRsNL8-CsVFCs-IHR0ClCF8
R
SWa)Q m_v7R 4:HRL0C_POs0FRR:=""jj;R--jRj:MlFsNlDRF;8CR:j4RHIs00C-EksFolERF;8CR:4jRNsC8C-LVCFs-HIs0lCRF
8C
RRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
R
RR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;1--Y,hBRYq1h
B
ShRQQ)a_qjv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_jRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_cRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_URR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_BRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
ShRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRR
R
RRRR2
;
RRRRuam)R
5
SmR7qm,7ARR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2O:=F_MP#_08DHFoOC_POs0F54j,U
2;
BSRp,iqBApi, RBq ,BAB,m mq,B, A)  1a)q, a1 A),W Wq,)R A:MRHR8#0_oDFH
O;
qSR7qq,7:ARRRHM#_08DHFoOC_POs0F5R4d8MFI0jFR2
;
SQR7qRR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;R

RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;S

RA7QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R
j2
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRX7ugRR:BbFlFMMC0#RHRk0sC
;









-
----------------------mb)v----------------------------B

mmvuha hRmb)v
R
RRRRt  h)RQB5
R
SRRRRaAQ_7WQa:]RR0HMCsoCR4:=;
S
SRRRRq) 7m_v7: RR0LHRR:=';j'
R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1h
B
SRRRRQQhaq_)vj_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R44:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R46:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R47:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.g:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vj_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd4:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_dRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vc_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd6:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_(RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vU_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdg:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ARR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vB_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd7:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_wRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RRRRRRRRR

R2RR;R

RuRRmR)a5S

RRRR7:mRR0FkR8#0_oDFHPO_CFO0s45dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;.2
R
SRBRRpRi,BR ,m,B R1)  :aRRRHM#_08DHFoO
;
SRRRRRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVbv)mRB:RFFlbM0CMRRH#0Csk;



----------------------------b--)Xmvg-R------------------------------------------
--
vBmu mhhbaR)Xmvg
R
RRRRt  h)RQB5
R
RRRRRRRRA_QaWaQ7]RR:HCM0oRCs:;=g
R
RRRRRR R)qv7_mR7 :HRL0=R:';j'
R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"R1--Y,hBRYq1h
B
RRRRRRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRR



RRRR
2;
RRRR)uma
R5
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2
;
SRRRRiBp, RB,BRm ),R a1 RH:RM0R#8F_Do;HO
R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV)RbmgvXRB:RFFlbM0CMRRH#0Csk;







-----------------------)-mv-------------------------
--
B

mmvuha hRv)mRR

RtRR )h Q5BRRS

RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SS

RRRR)7 q_7vm RR:LRH0:'=Rj
';
RRRRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YB-";-h1YBq,R1BYh
R
SRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRR
RR
RRRR
2;
RRRR)uma
R5
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsj.,d2
;
SRRRRiBp, RB, mB,1)  Wa,): RRRHM#_08DHFoO
;
RRRRSiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2
;
SRRRRRq7:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV)Rmv:FRBlMbFCRM0H0#Rs;kC




-
-----------------------------)Xmvg--------------------------------------------
-

m
Bvhum Rha)Xmvg
R
RRRRt  h)RQB5
R
RRRRRRRRA_QaWaQ7]RR:HCM0oRCs:;=g
R
RRRRRR R)qv7_mR7 :HRL0=R:';j'
R
RRRRRRpRAi _1pRR:L_H0P0COF:sR=jR"j;j"
R
RRRRRR R)1_ av m7R#:R0MsHo=R:RY"1h;B"-Y-1hRB,qh1YBR

RRRRRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRR



RRRR2
;
RRRRuam)R
5
SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd86RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsjn,d2
;
SpRBiB,R B,m  ,)1, aWR) :MRHR8#0_oDFH
O;
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;
qSR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVmR)vRXg:FRBlMbFCRM0H0#Rs;kC







---------------------------------1-s7-u--------------------------------------B

mmvuha hR7s1u
R
RRRRt  h)RQB5
R
SQRAaQ_W7_a]jRR:HCM0oRCs:n=4;R--4.,R,,RcRRU,4Rn,d
.
SQRAaQ_W7_a]4RR:HCM0oRCs:n=4;R--4.,R,,RcRRU,4Rn,d
.
S R)qv7_mR7 :HRL0=R:R''j;R--jL:R$#bN#FRl8RC;4b:RHDbCHRMClCF8
R
RRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R

RRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;-1BYh,1RqY
hB
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RR
R
RRRR2
;
RRRRuam)R
5
SmR7RF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsj.,d2
;
SpRBiBq,p,iARqB ,AB , mB,1)  ,aq)  1a:ARRRHM#_08DHFoO
;
S7Rqq7,qARR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj;R

RRRRA1pi :pRRRHM#_08DHFoOC_POs0F58.RF0IMF2Rj;S

RR7Q:MRHR8#0_oDFHPO_CFO0s45dRI8FMR0Fj
2
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVsu17RB:RFFlbM0CMRRH#0Csk;







--------------------------------s--1X7ug---------------------------------------
m
Bvhum Rhasu17X
gR
RRRRht  B)QR
5R
ASRQWa_Q]7a_:jRR0HMCsoCR4:=U-;-RRg,4RU,d
n
SQRAaQ_W7_a]4RR:HCM0oRCs:U=4;R--g4,RUd,RnS

Rq) 7m_v7: RR0LHRR:=';j'-j-R:$RLb#N#R8lFC4;R:HRbbHCDMlCRF
8C
ASRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R

RRRR)  1am_v7: RRs#0HRMo:"=R1BYh"-;-1BYh,1RqY
hB
QSRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvj:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv4:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qv.:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:.RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:dRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:nRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:(RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:qRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:ARR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd: RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
QSRh_Qa)_qvd:wRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjR"RRRRR
R
RR;R2
R
RRmRu)5aR
R
S7:mRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj=2:OPFM_8#0_oDFHPO_CFO0s,5jd;n2
R
SBqpi,iBpAB,R Bq, mA,B) , a1 q ,)1A aRH:RM0R#8F_Do;HO
R
Sq,7qqR7A:MRHR8#0_oDFHPO_CFO0sd54RI8FMR0Fj
2;
RRRRpRAip1 RH:RM0R#8F_Do_HOP0COF.s5RI8FMR0Fj
2;
7SRQRR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV1Rs7guXRB:RFFlbM0CMRRH#0Csk;







-----------------------sv)m----------------------------
m
Bvhum Rhasv)mRR

RtRR )h Q5BRRS

RRRRA_QaWaQ7]RR:HCM0oRCs:;=4SS

RRRR)7 q_7vm RR:LRH0:'=Rj
';
RRRRRRRRiAp_p1 RL:RHP0_CFO0s=R:Rj"jj
";
RRRRRRRR1)  va_mR7 :0R#soHMRR:="h1YB-";-h1YBq,R1BYh
R
SRQRRh_Qa)_qvj:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rj(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.d:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.A:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.w:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:jRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_4RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v._dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdd:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:cRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_6RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vn_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rd(:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:URR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_gRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vq_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdA:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:BRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_7RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v _dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdw:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"RRRRR
RR
RRRR
2;
RRRR)uma
R5
RSRRmR7RF:Rk#0R0D8_FOoH_OPC05Fsd84RF0IMF2Rj:F=OM#P_0D8_FOoH_OPC05Fsj.,d2
;
SRRRRiBp, RB,BRm ),R a1 RH:RM0R#8F_Do;HO
R
RRARSp i1pRR:H#MR0D8_FOoH_OPC05Fs.FR8IFM0R;j2
R
SRqRR7RR:H#MR0D8_FOoH_OPC05Fs48dRF0IMF2Rj
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRV)Rsm:vRRlBFbCFMMH0R#sR0k
C;




-

-----------------------------ms)v-Xg--------------------------------------------
m
Bvhum Rhasv)mX
gR
RRRRht  B)QR
5R
RRRRRRRRaAQ_7WQa:]RR0HMCsoCRg:=;R

RRRRR)RR _q7v m7RL:RH:0R=''j;R

RRRRRARRp1i_ :pRR0LH_OPC0RFs:"=Rj"jj;R

RRRRR)RR a1 _7vm RR:#H0sM:oR=1R"Y"hB;1--Y,hBRYq1h
B
RRRRRRRRQahQ_v)q_Rjj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rjc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RjB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvj:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qjv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_jRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R4B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv4:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q4v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_4RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.j:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.c:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.U:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_R.B:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qv.:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_q.v_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_.RL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdj:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:4RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_.RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vd_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_Rdc:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:6RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_nRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)v(_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdU:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:gRR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_qRR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vA_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj;S

RRRRQahQ_v)q_RdB:HRL0C_POs0FRR:=Xj"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj;j"
R
SRQRRh_Qa)_qvd:7RR0LH_OPC0RFs:X=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj
";
RSRRhRQQ)a_qdv_ RR:L_H0P0COF:sR="RXjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"
;
SRRRRQQhaq_)vw_dRL:RHP0_CFO0s=R:RjX"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjRRRRR



RRRR
2;
RRRR)uma
R5
7SRmRR:FRk0#_08DHFoOC_POs0F5Rd68MFI0jFR2O:=F_MP#_08DHFoOC_POs0F5dj,n
2;
BSRpRi,BR ,m,B R1)  :aRRRHM#_08DHFoO
;
RRRRRiAp1R p:MRHR8#0_oDFHPO_CFO0sR5.8MFI0jFR2
;
S7RqRH:RM0R#8F_Do_HOP0COF4s5dFR8IFM0R
j2
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRms)vRXg:FRBlMbFCRM0H0#Rs;kC








-
--------------------------q-u7U74-------------------------------------
--
vBmu mhhuaRq477US

SMoCCOsH5S

SRRRR q)tRR:LRH0:'=Rj-';-jR''L:R$#bN#FRl8RC;':4'RosCHC#0sRC8lCF8
S
SRRRRAt) RL:RH:0R=jR''
;R
RSSR1RRmt) RL:RH:0R=jR''
;
SRSRR7Rq7z_1ARR:LRH0:'=Rj
';
RRRRRRRRRRRR7uq7 _)1_ av m7R#:R0MsHo=R:RY"1h;B"-1-RY,hBqh1YBR

RRRRRRRRRARR1_ pv m7RL:RH:0R=4R''R--":4"RH#EVR0,":j"RsbNNCDDDMRHbRk0A
3
SRRRR
2;
RRRRRRR
R
RRRRRRFRbs
05
RSSRqRRRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SRRRRARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S

SRRRR q1pRR:H#MR0D8_FOoH;S

SRRRR,B B,pi)  1aRR:H#MR0D8_FOoH;S

SRRRR,1Q1RAQ:MRHR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;
RSSR1RRmA,1mRR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2
;
SRSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2
RRRRS
2;
7 hRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR7uq7R4U:FRBlMbFCRM0H0#Rs;kC







----------------------------u7q7g---------------------------------------
m
Bvhum Rhau7q7gR

RRRRRoRRCsMCH
O5
RSSRqRR)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8
C
SRSRR)RA :tRR0LHRR:=';j'RS

SRRRR)1m :tRR0LHRR:=';j'
S
SRRRRq_771RzA:HRL0=R:R''j;R

RRRRRRRRRuRRq_77)  1am_v7: RRs#0HRMo:"=R1BYh"-;-Rh1YB1,qY
hB
RRRRRRRRRRRR A1pm_v7: RR0LHRR:='-4'-4R""#:RE0HV,jR""b:RNDsNDRCDHkMb03RA
R
SR2RR;R

RRRRR
RR
RRRRFSbs50R
S
SRRRRqRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
S
SRRRRARR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
S
SRRRRqp1 RH:RM0R#8F_Do;HO
S
SRRRRBB ,p)i, a1 RH:RM0R#8F_Do;HO
S
SRRRR11Q,A:QRRRHM#_08DHFoOC_POs0F58URF0IMF2Rj;S

SRRRR,1m1RAm:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2;
RSSR7RRmRza:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2
SRRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFR7uq7:gRRlBFbCFMMH0R#sR0k
C;




-

-------------------------v--zgpaX-g----------------------------------
--
vBmu mhhvaRzgpaX
g
SCSoMHCsO
5
SRSRR)Rq :tRRHRL0=R:R''j;R--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8C
RSSRARR)R t:LRRH:0R=jR''
;
SRSRRzRma _)tRR:R0LHRR:=';j'
S
SRRRRu Qu_t) RR:RLRH0:'=Rj
';
RSSRqRR1hQt_t) RR:RLRH0:'=Rj
';
RSSRARR1hQt_t) RR:RLRH0:'=Rj
';
RRRRRRRRRRRRq1m_t) RR:RLRH0:'=RjR';
S
SRRRRvazp_1)  va_mR7 :0R#soHMRR:="h1YB-"-Rh1YBq,R1BYh
R
SR2RR;



RRRRFSbs50R
S
SRRRRqQ,1qRR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
S
SRRRRAQ,1ARR:H#MR0D8_FOoH_OPC05FsUFR8IFM0R;j2
S
SRRRRqt1QhA,R1hQtRH:RM0R#8F_Do;HO
R
RRRRRRRRRR1Rq Ap,1R p:MRHR8#0_oDFH
O;
RSSRBRR RR:H#MR0D8_FOoH;S

SRRRRiBpRH:RM0R#8F_Do;HO
S
SRRRR)  1aRR:H#MR0D8_FOoH;S

SRRRRz7maRR:FRk0#_08DHFoOC_POs0F5R4(8MFI0jFR2
;
RRRRRRRRRRRR1,mq1RmA:kRF00R#8F_Do_HOP0COFUs5RI8FMR0Fj
2
SRRRR
2;
7 hRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvzaggXRB:RFFlbM0CMRRH#0Csk;







----------------------------pvzaX4U4-U--------------------------------------



vBmu mhhvaRz4paUUX4
R
RRCRoMHCsO
5
S)Sq :tRRHRL0=R:R''j;R--R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8C
ASS)R t:LRRH:0R=jR''
;
SzSma _)tRR:R0LHRR:=';j'
S
Su Qu_t) RR:RLRH0:'=Rj
';
qSS1hQt_t) RR:RLRH0:'=Rj
';
ASS1hQt_t) RR:RLRH0:'=Rj
';
RRRRRRRRq1m_t) RR:RLRH0:'=Rj
';
vSSz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"R--1BYh,1RqY
hB
;S2



SsbF0
R5
qSS,q1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SAQ,1ARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S

SQq1tRh,At1QhRR:H#MR0D8_FOoH;R

RRRRRqRR1, pAp1 RH:RM0R#8F_Do;HO
S
SB: RRRHM#_08DHFoO
;
SpSBiRR:H#MR0D8_FOoH;S

S1)  :aRRRHM#_08DHFoO
;
SmS7z:aRR0FkR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;
RRRRRRRRq1m,A1mRF:Rk#0R0D8_FOoH_OPC05Fs48(RF0IMF2Rj
2
S;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFvVRz4paUUX4RB:RFFlbM0CMRRH#0Csk;







----------------------------pvzaXdnd-n--------------------------------------B

mmvuha hRpvzaXdnd
n
SMoCCOsH5S

S q)tRR:R0LHRR:=';j'-R-R':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8
C
S)SA :tRRHRL0=R:R''j;S

Samzj _)tRR:R0LHRR:=';j'
S
Sm4za_t) RR:RLRH0:'=Rj
';
uSSQ_u )R t:LRRH:0R=jR''
;
S1SqQ_th)R t:LRRH:0R=jR''
;
S1SAQ_th)R t:LRRH:0R=jR''
;
SzSvp)a_ a1 _7vm RR:#H0sM:oR=1R"Y"hB-1-RY,hBRYq1h
B
S
2;
S

b0FsR
5
SRSq:MRHR8#0_oDFHPO_CFO0s65dRI8FMR0Fj
2;
ASSRH:RM0R#8F_Do_HOP0COFds56FR8IFM0R;j2
S
Sqt1QhA,R1hQtRH:RM0R#8F_Do;HO
S
SB: RRRHM#_08DHFoO
;
SpSBiRR:H#MR0D8_FOoH;S

S1)  :aRRRHM#_08DHFoO
;
SmS7z:aRR0FkR8#0_oDFHPO_CFO0s45(RI8FMR0Fj
2
S
2;
7 hRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvzaXdnd:nRRlBFbCFMMH0R#sR0k
C;




-

-------------------------v--zqpapnzdX-4U-------------------------------------
-
Bumvmhh azRvppaqzXdn4
U
SMoCCOsH5S

S q)tRR:R0LHRR:=';j'-R-R':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8
C
S)SA :tRRHRL0=R:R''j;S

S B)tRR:R0LHRR:=';j'
S
Sm_za)R t:LRRH:0R=jR''
;
SQSuu) _ :tRRHRL0=R:R''j;S

SQq1t)h_ :tRRHRL0=R:R''j;S

SQA1t)h_ :tRRHRL0=R:R''j;R

RRRRRqRRBmBpq)7_ Rtj:HRL0=R:R''j;R

RRRRRqRRBmBpq)7_ Rt4:HRL0=R:R''j;R

RRRRR1RRm)q_ :tRR0LHRR:=';j'
R
RRRRRRzRvppaqzXdn4vU_mR7 :MRH0CCos=R:R-j;-dj:nUG4R-+/RRB;4B:qBR/j+nRdG;4URR.:d4nGURR+BQq1
R
RRRRRR_RBq_771RzA:HRL0=R:R''j;R--':j'R8N8;'RR4R':#
kL
vSSz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"R--1BYh,1RqY
hB
;S2
R
RR
R
SsbF0
R5
qSSRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SARR:H#MR0D8_FOoH_OPC05Fsd86RF0IMF2Rj;S

S:BRRRHM#_08DHFoOC_POs0F5R6d8MFI0jFR2
;
S1SqQ,thRQA1tRh,qpBBmRq7:MRHR8#0_oDFH
O;
BSS RR:H#MR0D8_FOoH;S

SiBpRH:RM0R#8F_Do;HO
S
S)  1aRR:H#MR0D8_FOoH;S

S1BqQRR:H#MR0D8_FOoH_OPC05Fs68cRF0IMF2Rj;S

Sz7maRR:FRk0#_08DHFoOC_POs0F5R6d8MFI0jFR2
;
SqSB1:mRR0FkR8#0_oDFHPO_CFO0sc56RI8FMR0Fj
2
S
2;
7 hRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRpvzazqpd4nXURR:BbFlFMMC0#RHRk0sC
;
RRRR




-
--------------------------z-vp7aq7zqp44UXU---------------------------------------
m
Bvhum Rhavazpqq77pUz4X
4U
CSoMHCsO
5
SjSq)R t:HRL0=R:R''j;R--':j'RbL$NR##lCF8;4R''s:RC#oH0CCs8FRl8
C
SjSA)R t:HRL0=R:R''j;
R
S4Sq)R t:HRL0=R:R''j;S

S)A4 :tRR0LHRR:=';j'
S
SBt) RL:RH:0R=jR''
;
SzSma _)tRR:LRH0:'=Rj
';
uSSQju _t) RL:RH:0R=jR''
;
SQSuu_ 4)R t:HRL0=R:R''j;S

SQq1t_hj)R t:HRL0=R:R''j;S

SQA1t_hj)R t:HRL0=R:R''j;S

SQq1t_h4)R t:HRL0=R:R''j;S

SQA1t_h4)R t:HRL0=R:R''j;S

SBqBp7mq_t) jRR:LRH0:'=Rj
';
qSSBmBpq)7_ Rt4:HRL0=R:R''j;R

RRRRR1RRm)q_ :tRR0LHRR:=';j'
S
SA7_q7z_1ARR:LRH0:'=Rj-';-jR''N:R8R8;':4'RL#k
S
SB7_q7z_1ARR:LRH0:'=Rj
';
vSSzqpa7p7qzX4U4vU_mR7 :MRH0CCos=R:R-j;-4j:UUG4R-+/RG4U4+UR/B-R;4RR:BRqBR/j+UR4GR4U+R/-44UGU.;R:G4U4+UR/4-RUUG4RB+Rq
1Q
vSSz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"R--1BYh,1RqY
hB
;S2



SsbF0
R5
qSSj4,qRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SAAj,4RR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S

Sq1Q,A1QRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SBRR:H#MR0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R

RRRRRqRR1hQt,QA1t:hRRRHM#_08DHFoOC_POs0F584RF0IMF2Rj;R

RRRRRqRR1, pAp1 RH:RM0R#8F_Do_HOP0COF4s5RI8FMR0Fj
2;
RRRRRRRR1BqQRR:H#MR0D8_FOoH_OPC05Fs68cRF0IMF2Rj;R

RRRRRqRRBmBpq:7RRRHM#_08DHFoO
;
S SBRH:RM0R#8F_Do;HO
S
SBRpi:MRHR8#0_oDFH
O;
)SS a1 RH:RM0R#8F_Do;HO
S
S7amzRF:Rk#0R0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R

RRRRR1RRm1q,m:ARR0FkR8#0_oDFHPO_CFO0s(54RI8FMR0Fj
2;
BSSqR1m:kRF00R#8F_Do_HOP0COF6s5cFR8IFM0R
j2
;S2
h
 7mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvp7aq7zqp44UXURR:BbFlFMMC0#RHRk0sC
;





-
--------------------------z-vppaqzX4U4-U--------------------------------------B

mmvuha hRpvzazqp44UXUS

oCCMs5HO
S
Sqt) RL:RH:0R=jR''-;-R''j:$RLb#N#R8lFC';R4R':sHCo#s0CCl8RF
8C
ASS)R t:HRL0=R:R''j;
R
S)SB :tRR0LHRR:=';j'
S
S7t) RL:RH:0R=jR''
;
RRRRRRRRm_za)R t:HRL0=R:R''j;S

SuuQ  _)tRR:LRH0:'=Rj
';
qSS1hQt_t) RL:RH:0R=jR''
;
S1SAQ_th)R t:HRL0=R:R''j;S

SQ71t)h_ :tRR0LHRR:=';j'
S
SqpBBm_q7)j tRL:RH:0R=jR''
;
SBSqBqpm7 _)t:4RR0LHRR:=';j'
S
SA7_q7z_1ARR:LRH0:'=Rj-';-jR''N:R8R8;':4'RL#k
S
SB7_q7z_1ARR:LRH0:'=Rj
';
vSSzqpapUz4X_4Uv m7RH:RMo0CC:sR=;Rj-:-jq/BBj/R+-UR4GR4U+R/-B4;R:BqB/+jR/4-RUUG4RB+Rq;1QRR.:44UGU/R+-RR7+qRB1
Q;
vSSz_pa)  1am_v7: RRs#0HRMo:"=R1BYh"R--1BYh,1RqY
hB
;S2



SsbF0
R5
qSSRH:RM0R#8F_Do_HOP0COF4s5(FR8IFM0R;j2
S
SARR:H#MR0D8_FOoH_OPC05Fs48(RF0IMF2Rj;S

SRB,7RR:H#MR0D8_FOoH_OPC05Fs68dRF0IMF2Rj;R

RRRRRqRR1hQt,1RAQRth:MRHR8#0_oDFH
O;
RRRRRRRR1BqQRR:H#MR0D8_FOoH_OPC05Fs68cRF0IMF2Rj;R

RRRRRqRRBmBpq77,1hQtRH:RM0R#8F_Do;HO
S
SB: RRRHM#_08DHFoO
;
SpSBiRR:H#MR0D8_FOoH;S

S1)  :aRRRHM#_08DHFoO
;
SmS7z:aRR0FkR8#0_oDFHPO_CFO0sd56RI8FMR0Fj
2;
BSSqR1m:kRF00R#8F_Do_HOP0COF6s5cFR8IFM0R
j2
;S2
h
 7mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVzRvppaqzX4U4:URRlBFbCFMMH0R#sR0k
C;




-

-------------------------q--pcz67------------------------------------
--
vBmu mhhqaRpcz67S

oCCMs5HO
R
SRqRR)R t:HRL0=R:R''j;'--jR':LN$b#l#RF;8CR''4:CRso0H#C8sCR8lFCR

RRRRRARR)R t:HRL0=R:R''j;S

RRRRqt1Qh _)tRR:LRH0:'=Rj
';
RSRR1RAQ_th)R t:HRL0=R:R''j;S

RRRRqpBBm_q7)R t:HRL0=R:R''j;S

RRRRm_za)R t:HRL0=R:R''j;S

RRRRA7_q7z_1ARR:LRH0:'=Rj-';-''j:8N8;4R''k:#LS

RRRRB7_q7z_1ARR:LRH0:'=Rj
';
RRRRRRRRzqp7m_v7: RR0HMCsoCRR:=j-;-jB:qBR/j+R/-A/R+-;RqRq4:BjB/R-+/R+ARR1BqQ.;R:+qR/A-RRB+Rq;1Q
S
Sq_pz)  1am_v7: RRs#0HRMo:"=R1BYh"1--Y,hBRYq1h
B
RRRR2
;
RRRRb0FsR
5
SRRRR:qRRRHM#_08DHFoOC_POs0FRd56RI8FMR0Fj
2;
RSRRRRA:MRHR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
R
SRBRR RR:H#MR0D8_FOoH;S

RRRRBRpi:MRHR8#0_oDFH
O;
RSRR R)1R a:MRHR8#0_oDFH
O;
RSRR1RqQ,thAt1QhRR:H#MR0D8_FOoH;S

RRRRqpBBmRq7:MRHR8#0_oDFH
O;
RSRRqRB1:QRRRHM#_08DHFoOC_POs0FRc56RI8FMR0Fj
2;
RSRRmR7z:aRR0FkR8#0_oDFHPO_CFO0s6R5dFR8IFM0R;j2
R
SRBRRqR1m:kRF00R#8F_Do_HOP0COF5sR68cRF0IMF2Rj
R
RR;R2
h
 7mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRqz76cRB:RFFlbM0CMRRH#0Csk;







--------------------z-Aw-t--------------------------



vBmu mhhAaRzRwt
R
Ruam)5R

RSRRmRR:FRk0#_08DHFoO
;
RRRRS:QRRRHM#_08DHFoOR

R2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGFAVRzRwt:FRBlMbFCRM0H0#Rs;kC




-
--------------A--z-w1-----------------
--
B

mmvuha hRwAz1
R
RRRRuam)R
5
RRRRRRRRR:mRR0FkR8#0_oDFH
O;
RRRRRRRRRRQ:MRHR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVA1zwRB:RFFlbM0CMRRH#0Csk;



-

---------------------7th-----------------



vBmu mhhtaRh
7R
RRRR)uma
R5
RRRRtSRRF:Rk#0R0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVhRt7RR:BbFlFMMC0#RHRk0sC
;




---------------------BeB------------------------



Bumvmhh aBReB
R
RRRRuam)R
5
RRRRSRRe:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRBeBRB:RFFlbM0CMRRH#0Csk;







----------------------------t--1-)--------------------------------------



vBmu mhhtaR1
)R
RRRR)uma
R5
RRRRRRRR1Rt):QRRRHM#_08DHFoOR

R2RR;C

MB8Rmmvuha h;



0SN0LsHkR0C#_$MLODN	F_LGVRFR)t1RB:RFFlbM0CMRRH#0Csk;R

RNRR0H0sLCk0RM#$_bMFsCkMRRFVtR1):FRBlMbFCRM0H0#Rs;kC




-
-----------------m-1B-------------------------
--
vBmu mhhmaR1
BR
RRRRht  B)QR
5
RRRRRRRRwT) _e7QRH:RMo0CC:sR=jR4j-;-..~4UM,FDC$RPRCMM
kl
RRRRRRRRe7 QRB :0R#soHMRR:="4tWh"-.-W-t4.h-,4tWh,-cthW4-tn,W-4hgW,t4-h)cW,t4-h)gW,t4.h-AW,t4ch-AW,t4-h)ctA,W-4hn, 1thW4-1g ,4tWhg)- 
1
RRRR2
;
RRRRuam)R
5
SRRRRBm1mRza:kRF00R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRBm1RB:RFFlbM0CMRRH#0Csk;







--------------------------------pup-------------------------
-
Bumvmhh apRupR

RtRR )h Q
B5
RRRRRRRRRRRRBRwphiQR1:Rah)Qt=R:Rj"4j"3j;V--skCJC$MORRFV0RECOHD	M25v
R
RRRRRRRRRR7RR BeQ RR:1Qa)h:tR=tR"W-4h.-";-W"t44h-"t,"W-4h."",thW4-,c""4tWh"-n,tR"W-4hg"",thW4)"-c,W"t4-h)g"",thW4-".A,W"t4ch-A"",thW4)A-c"t,"W-4hn" 1,W"t4gh- ,1""4tWhg)- ,1""4tWh.1-"t,"W14h-".B,W"t4-hZ4"",thW41.)-B"",thW4-"41,W"t4 h1-".B
R
RRRRRRRRRR7RRYQh_7_Qe1R p:aR1)tQhRR:="DVN#;C"-s-0kQC:7p1 ;NRVD:#CQe7Q_p1 
R
RRRRRRRRRRQRR7_Qe1R p:MRH0CCos=R:R-j;-bQMk80RH8PHCQsR7,QeR4j:,.4:3n33dc:n34RR~
nc
RRRRRRRRRRRRYR7hA_w7_Qe1R p:aR1)tQhRR:="DVN#;C"
R
RRRRRRRRRRwRRAe7Q_p1 RH:RMo0CC:sR=;Rj-C-wCN8LO8	RH8PHCwsRAe7Q,jRR:44,:3.33:ndnRc34c~n
R
RRRRRRRRRR7RRYmh_7_Qe1R p:aR1)tQhRR:="DVN#;C"-s-0kmC:7p1 ;NRVD:#Cme7Q_p1 
R
RRRRRRRRRRmRR7_Qe1R p:MRH0CCos=R:R-U;-c.//4U/n./d//cUnUc/jn/g/.44/U4.
R
RRRRRRRRRRuRR1_7q1R p:aR1)tQhRR:="jjjj-";-R

RRRRRRRRRRRR7_Yh7 q_hRR:1Qa)h:tR=VR"NCD#"-;-0Csk:7u1qsRFRa7zYR7qFwsR7Rq;V#NDC7:Rq _1pR

RRRRRRRRRRRR7Yza71q_ :pRR)1aQRht:"=R4jjj"-;-
R
RRRRRRRRRRBRRpzimaa_w_)7QRL:RH:0R=4R''-;-RiBpmRzaVCHMRM0kHRMo8CHsOF0HM'3R4F'RMRD$
R
RRRRRRRRRRBRRpzimawu_aQ_7)RR:LRH0:'=R4-';-4R''MRFD
$
RRRRRRRRRRRRRiBpm_za7_pY1ua RH:RMo0CC:sR=;Rj-j-R,.4,,
c
RRRRRRRRRRRRRiBpmuza_Y7p_ 1auRR:HCM0oRCs:j=R;R--j,,4.



RRRRRRRRRRRRpRBiamz71d_):BRR)1aQRht:"=RBmpiz;a"-C-#D0CORP8HdkRF00bk,pRBiamzusRFRiBpm
za
RRRRRRRRRRRRpRBi_wA1R p:aR1)tQhRR:="0HMCNsMD
";
RRRRRRRRRRRRpRBiamz_uAYqR11:aR1)tQhRR:="DVN#;C"
R
RRRRRRRRRRBRRpzimaAu_Y1uq1RR:1Qa)h:tR=VR"NCD#"
;
RRRRRRRRRRRRRiBpm7za_uAYqR11:aR1)tQhRR:="DVN#;C"
R
RRRRRRRRRRBRRpzima17_):BRR)1aQRht:"=RBmpiz;a"-C-#D0CORP8HR0Fkb,k0RpRBiamzusRFRiBpm
za
RRRRRRRRRRRRYR7h7_1Q1e_ :pRR0HMCsoCRR:=.R--..~4UM,FDC$RPRCMM
kl
RRRRRRRRRRRR
R
SRRRR2RR;R

RuRRm5)a
R
RRRRRRRRRRBRRphiQRQ:Rh0R#8F_Do;HO
R
RRRRRRRRRRBRRpAiwRQ:Rh0R#8F_Do:HO=''j;R

RRRRRRRRRRRRQ 71pRR:Q#MR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
R
RRRRRRRRRRwRRA 71pRR:Q#MR0D8_FOoH_OPC05Fs6FR8IFM0R;j2
R
RRRRRRRRRRmRR7p1 RQ:RM0R#8F_Do_HOP0COF6s5RI8FMR0Fj
2;
RRRRRRRRRRRR R)1R a:MRHR8#0_oDFH=O:';j'
R
RRRRRRRRRR)RR a1 _:uRRRHM#_08DHFoO':=j
';
RRRRRRRRRRRR R)1_ aQHR:M0R#8F_Do:HO=''j;R

RRRRRRRRRRRR)  1aR_1:MRHR8#0_oDFH:OR=''j;R

RRRRRRRRRRRRuq17,pw7YRR:Q#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
R
RRRRRRRRRR7RRz7aYqRR:Q#MR0D8_FOoH_OPC05FsdFR8IFM0R;j2
R
RRRRRRRRRRpRRmRBi:zRma0R#8F_Do;HO
R
RRRRRRRRRRBRRpzimaRR:mRza#_08DHFoO
;
RRRRRRRRRRRRRiBpm7zaRF:Rk#0R0D8_FOoH;R

RRRRRRRRRRRRBmpizRau:kRF00R#8F_Do;HO
R
RRRRRRRRRRBRRpzimaR7d:kRF00R#8F_Do
HO
RRRRRRRR
2;
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRpupRB:RFFlbM0CMRRH#0Csk;







----------------p-ae_71QwAz---------------------------------



vBmu mhhaaRp1e7_zQAwR

RuRRm5)a
R
RRRRRRRRm:zRma0R#8F_Do;HO
R
RRRRRRRRQ:hRQR8#0_oDFH
O;
RRRRRRRRRQA:hRQR8#0_oDFH
O
RRRRRRRR2
;
CRM8Bumvmhh a
;
RRRRNs00H0LkC$R#MD_LN_O	LRFGFaVRp1e7_zQAwRR:BbFlFMMC0#RHRk0sC
;
RRRRNs00H0LkCDRLN_O	L_FGb_N8bRHMFaVRp1e7_zQAwRR:BbFlFMMC0#RHR,"QR"QA;







----------------p-ae_71mwAz---------------------------------



vBmu mhhaaRp1e7_zmAwR

RuRRm5)a
R
RRRRRRRRm:zRma0R#8F_Do;HO
R
RRRRRRARmRm:Rz#aR0D8_FOoH;R

RRRRRQRRRQ:Rh0R#8F_Do
HO
RRRRRRRR
2;
8CMRvBmu mhh
a;
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFVa7pe1A_mz:wRRlBFbCFMMH0R#sR0k
C;
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFVa7pe1A_mz:wRRlBFbCFMMH0R#mR",ARm"
;





-
--------------a--p1e7_zaAw--------------------------------
-

m
Bvhum Rhaa7pe1A_az
w
RRRRuam)R
5
RRRRSRRmRm:RzRaRR8#0_oDFH
O;
RRRRmSRARR:mRza#_08DHFoO
;
RRRRRQSRRRR:QRhRR0R#8F_Do;HO
R
SRRRRmR h:hRQRRRR#_08DHFoOR

R2RR;C

MB8Rmmvuha h;R

RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpRae_71awAzRB:RFFlbM0CMRRH#0Csk;R

RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpRae_71awAzRB:RFFlbM0CMRRH#"Rm,m;A"







-----------------eap7Q1_mwAz---------------------------------



vBmu mhhaaRp1e7_AQmz
w
RRRRuam)R
5
RRRRSRRmRm:RzRaRR8#0_oDFH
O;
RRRRQSRm:ARRmQhz#aR0D8_FOoH;R

RRRRRRRRQ:mRRmQhz#aR0D8_FOoH;R

RRRRSRRQRQ:RhRRRR8#0_oDFH
O;
RSRRmRR :hRRRQhR#RR0D8_FOoH
R
RR;R2
M
C8mRBvhum ;ha
R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFReap7Q1_mwAzRB:RFFlbM0CMRRH#0Csk;R

RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpRae_71QzmAwRR:BbFlFMMC0#RHRm"Q,mRQA
";




-

---------------- 7pe1A_Qz-w------------------------------
--
B

mmvuha hRe p7Q1_A
zw
RRRR)uma
5
RRRRRRRRmRR:mRza#_08DHFoO
;
RRRRRRRRQRR:Q#hR0D8_FOoH;R

RRRRRQRRARR:Q#hR0D8_FOoH
R
RRRRRR;R2
M
C8mRBvhum ;ha
R
RR0RN0LsHkR0C#_$MLODN	F_LGVRFRe p7Q1_ARzw:FRBlMbFCRM0H0#Rs;kC
R
RR0RN0LsHkR0CLODN	F_LGN_b8H_bMVRFRe p7Q1_ARzw:FRBlMbFCRM0H"#RQQ,RA
";




-

---------------- 7pe1A_mz-w------------------------------
--
B

mmvuha hRe p7m1_A
zw
RRRR)uma
5
RRRRRRRRmRR:mRza#_08DHFoO
;
RRRRRRRRm:ARRamzR8#0_oDFH
O;
RRRRRRRR:QRRRQh#_08DHFoOR

RRRRR2RR;C

MB8Rmmvuha h;R

RNRR0H0sLCk0RM#$_NLDOL	_FFGRVpR e_71mwAzRB:RFFlbM0CMRRH#0Csk;R

RNRR0H0sLCk0RNLDOL	_FbG_Nb8_HFMRVpR e_71mwAzRB:RFFlbM0CMRRH#"Rm,m;A"







-----------------e p7a1_A-zw--------------------------------



Bumvmhh apR e_71awAz
R
RRmRu)5aR
R
RRRRSm:RRRamzR#RR0D8_FOoH;R

RSRRRRmA:zRma0R#8F_Do;HO
R
RRSRRRRQR:hRQRRRR#_08DHFoO
;
SRRRR RmhRR:QRhRR0R#8F_Do
HO
RRRR
2;
8CMRvBmu mhh
a;
RRRR0N0skHL0#CR$LM_D	NO_GLFRRFV 7pe1A_az:wRRlBFbCFMMH0R#sR0k
C;
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1A_az:wRRlBFbCFMMH0R#mR",ARm"
;





-
-------------- --p1e7_AQmz-w------------------------------
--
B

mmvuha hRe p7Q1_mwAz
R
RRmRu)5aR
R
RRRRSm:RRRamzR#RR0D8_FOoH;R

RSRRRAQmRQ:RhamzR8#0_oDFH
O;
RRRRRRRRmRQRQ:RhamzR8#0_oDFH
O;
RRRRRRSQ:RRRRQhR#RR0D8_FOoH;S

RRRRRhm RQ:RhRRRR8#0_oDFH
O
RRRR2
;
CRM8Bumvmhh a
;
RRRRNs00H0LkC$R#MD_LN_O	LRFGF VRp1e7_AQmz:wRRlBFbCFMMH0R#sR0k
C;
RRRR0N0skHL0LCRD	NO_GLF_8bN_MbHRRFV 7pe1m_QARzw:FRBlMbFCRM0H"#RQRm,Q"mA;







--------------------------------iBp7-Qe-------------------------B

mmvuha hRiBp7
Qe
RRRRht  B)Q5S

RRRRRe7Q_7vm RR:1Qa)h:tR=.R""-;-R"".,dR"3,6"R""c,6R""",RU""5Um",MRD$#bkbFCs08MRHR4oIM	-n/,g	oMI4#	-.,4oIM#-42S

RRRRR)t1 :hRR)1aQRht:"=RV#NDC-"-RN"VD"#C,0R"s"kC
R
SR2RR;R

RuRRm5)a
R
RRRRRR]RRBQpihRR:Q#hR0D8_FOoH;S

RRRRR1)  Rah:hRQR8#0_oDFH
O;
RSRRBRRqApQRQ:RM0R#8F_Do;HO
R
SRRRRBmpiz:aRRamzR8#0_oDFH
O
RRRRRRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFVB7piQ:eRRlBFbCFMMH0R#sR0k
C;




-

----------------7-pp--------------------------------
m
Bvhum Rha7
pp
RRRRht  B)Q5R

RRRRR7RRpwp_m )BRH:RMo0CC:sR=;Rj-:-4RsVFODCRFRO	NRM8OCF8;:RjR8OFCF/DOo	RCsMCN80CRFVslpR7pFRDF
b
RRRRRRRR7_Qe1R p:HRL0=R:R''4;j--,sMFlRNDD	FOR8lFC4;R,#VN0FRDOl	RF
8C
RSRRmRB7B 1q:pRR)1aQRht:"=Rj"jj;j--jj4R4jjR444Rj4jRj44R44jR4
4
RRRRRRRR1pBq_R h:aR1)tQhRR:="k0sC-"-0Csk,DVN#
C
RRRR2
;
RRRRuam)5R

RRRRRBRRphiQ:RQh#_08DHFoO':=j
';
RRRRRRRRm1auQ:RM0R#8F_Do:HO=''j;R

RRRRR)RR a1 RQ:RM0R#8F_Do:HO=''j;R

RRRRRzRRuB7hhRap:MRQR8#0_oDFH=O:';j'
R
RRRRRRmRpB:iRRamzR8#0_oDFH
O;
RRRRRRRR 1auRR:mRza#_08DHFoOC_POs0F58(RF0IMF2Rj
R
RR2RR;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRp:pRRlBFbCFMMH0R#sR0k
C;




-

-----------------------------p7p7-pY-------------------------------------
-
Bumvmhh apR7pY7p
R
RR RthQ )B
5
RRRRRRRR7_ppQ h1pRR:LRH0:'=Rj-';-''j:bL$NR##lCF8,4R''k:R#8CRD8D_C$DNRDOCDR

RRRRR7RRp1Y_QRth:HRL0=R:R''j;R--':j'',+'R4R''':R-
'
RRRRRRRR7_pYqR7K:MRH0CCos=R:R-j-j6~.68,RD#$_H=oMj8R:DN$_8R[;8_D$#MHo=-4:.+6n8_D$N
8[
RRRR
2;
RRRR)uma
5
RRRRRRRR71ppaR u:hRQR8#0_oDFHPO_CFO0sR5(8MFI0jFR2
;
RRRRRRRRBQpihh:QR8#0_oDFH
O;
RRRRRRRR)7Q,qpm7vh,m:e RRQM#_08DHFoO
;
RRRRRRRRBmpiz:aRRamzR8#0_oDFH
O;
RRRRRRRRqwptRR:mRza#_08DHFoOR

RRRR2
;
CRM8Bumvmhh a
;
S0N0skHL0#CR$LM_D	NO_GLFRRFV77ppp:YRRlBFbCFMMH0R#sR0k
C;




-

-----------------------------qwp16].n-i--------------------------------------B

mmvuha hRqwp16].n
i
RRRRuam)5R

RRRRRXRRqR7):hRQR8#0_oDFHPO_CFO0sR5n8MFI0jFR2
;
RRRRRRRRY)q7RQ:Rh0R#8F_Do_HOP0COF6s5RI8FMR0Fj
2;
RRRRRRRR,X Y1 , h:QR8#0_oDFH
O;
RRRRRRRRh7QRQ:Rh0R#8F_Do_HOP0COFds54FR8IFM0R;j2
R
RRRRRR)R q,1 ut)m,1heaR):Q#hR0D8_FOoH;R

RRRRR7RRmRza:zRma0R#8F_Do_HOP0COFds54FR8IFM0R
j2
RRRR;R2
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVpRwq.1]6Rni:FRBlMbFCRM0H0#Rs;kCRRRR







--------------------------------7 ]Bh------------------------------------
-
Bumvmhh a]R7B
 h
RRRR)uma
R5
BSRpzimaRR:mRza#_08DHFoO
;S
BSR RR:Q#hR0D8_FOoH;
S
SpRBiRQh:hRQR8#0_oDFH
O
RRRR2
;S
8CMRvBmu mhh
a;
0SN0LsHkR0C#_$MLODN	F_LGVRFRB7] :hRRlBFbCFMMH0R#sR0kRC;R
RR




-

--------------------------------7-B1------------------------------------
m
Bvhum Rha7
B1
RRRRht  B)QR
5
SBS71m_v7: RRs#0HRMo:"=R)QQ1h-t"-iBpjp,BiB4,p,i.Bdpi,7th,BeB,1)QQ,htwpqpQ,htBjpi_7th,iBpjB_eBp,Bit4_hB7,p_i4e,BBB.pi_7th,iBp.B_eBp,Bitd_hB7,p_ide
BB
;S2
u
SmR)a5S

SiBpjRR:Q#hR0D8_FOoH;S

SiBp4RR:Q#hR0D8_FOoH;S

SiBp.RR:Q#hR0D8_FOoH;S

SiBpdRR:Q#hR0D8_FOoH;S

SiBp1R p:hRQR8#0_oDFHPO_CFO0sR5d8MFI0jFR2
;
S S1p)wmB: RRRQh#_08DHFoO
;
SpSBiamzRm:Rz#aR0D8_FOoH
2
S;C

MB8Rmmvuha h;S

Ns00H0LkC$R#MD_LN_O	LRFGF7VRB:1RRlBFbCFMMH0R#sR0kRC;R
RR




-

-----------------------------7--T-B ------------------------------------
m
Bvhum Rha7 TB
R
RRmRu)5aR
R
SBmpiz:aRRamzR8#0_oDFHSO;
R
SB: RRRQh#_08DHFoO
;S
BSRphiQRQ:Rh0R#8F_Do
HO
RRRRS2;
M
C8mRBvhum ;ha
N
S0H0sLCk0RM#$_NLDOL	_FFGRVTR7B: RRlBFbCFMMH0R#sR0kRC;R
RR




C

MB8Rmmvuha h1
;





