--=============================== entity and architecture dw_div===============================
@E-

-------------------------------------------------------------------------------------------------
-----
-HRa0RDCRRRRRRR:78W_H-P
-CR7#MHoRRRRRRR:78W_H-P
-kRq0sEFRRRRRRR:1PCDN)lRR]/RN#sHERRvi-
-RlBFb$NMRRRRR1:R$DMbH0OH$FR1VN0IsQCRMN8HR0uP30Rp8-3
--
---------------------------------------------------------------------------------------------------
-R#7CObsH0MHFR7:RWH_8P#RHRONRFHlLMHN0FDMNR0HMCsoCRP8HHs8CR0IHEFSL0JERkHF0CRM0NRM8sNClHCM8skRF00bk#
3R-a-RERH#ObFlFMMC0HR8PCH8#ER0CHR8PCH8MR8,NL,R$ER0CHR8PFH#sL,R,FR0RFbs8CkORC0ERFJk0MHC0MRN8CRslMNH83Cs
R--mHb0FDMNDR$,0RECsNClHCM8skRF00bkRlOFbCk0#ER0CFRl8kkD#-3
--
-RCaERo#HMVRFRC0ERlsCN8HMCHsR#ER0CHR#oFMRVER0CRRqHkMb0-3
-ERaCHR#oFMRVER0CFRl8kkD##RHRC0ERo#HMVRFRC0ERHARM0bk3-
-
R--)HCP#MHFR#]H0$Fs
R--j4c/(./4RC51DlPN2w:RH8GCRoDFHHOR#C#kRsVFR0LFEkRTFC0HMN0RM)8RCHlNMs8CRsVFRC0ER#ONCVRFRP8HHM8HoHRI0-ER4#R5HCoM8bRFC0sNH2FM
---------------------------------------------------------------------------------------------------


SDsHLNRs$Q   ;#
kC RQ # 30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;kR#CHCCC38#0_oDFHNO_sEH03DND;C

M00H$WR7_P8HR
H#SMoCCOsH5S
SNH_I8S0ERm:u1QQae: S=;4c
LSS_8IH0RES:1umQeaQ =S:gS;
S_0OlCF8ShR:q)azqSpR:;=j
sSSCll_FR8C:ahqzp)qS4:=
2SS;b
SF5s0
NSSRSSS:MRHR8#0_oDFHPO_CFO0s_5NI0H8ER-48MFI0jFR2S;
SSLRSRS:H#MR0D8_FOoH_OPC05FsLH_I8-0E4FR8IFM0R;j2
JSSkHF0CSM0:kRF00R#8F_Do_HOP0COFNs5_8IH04E-RI8FMR0Fj
2;SCSslMNH8SCs:kRF00R#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;SHS8PCH8__L$jRS:FRk0#_08DHFoOS
S2C;
M78RWH_8P
R;
ONsECH0Os0kC0RsDVRFR_7W8RHPH
#R
R--QCM0sDMNRo#HMRND8DCON0sNH#FM
o#HMRNDbNNslR4,J0kF,kRJFC0HM.0_#0,RCRlb:0R#8F_Do_HOP0COF5sRRIN_HE80R4-RRI8FMR0Fj;R2
o#HMRNDbNNslR.,lDF8R#:R0D8_FOoH_OPC0RFs5_RLI0H8ERR-4FR8IFM0R2jR;
R
-w-Rk0MOHRFM0oFRC00REJCRkHF0CRM0NRM8sNClHCM8s13RE0HV/L#k#N0sOM0RFsMRCF#0soHMRoNDF0sHEHlR#lRHblDCCCM08

SVOkM0MHFRP8HRN5RR#:R0D8_FOoH_OPC05FsRIN_HE80R4-RRI8FMR0Fj;R2R:LRR8#0_oDFHPO_CFO0sL5R_8IH0-ERR84RF0IMFRRj2RR2skC0s#MR0D8_FOoH_OPC0;Fs
k
VMHO0F8MRH5PRR:NRR8#0_oDFHPO_CFO0sN5R_8IH0-ERR84RF0IMFRRj2L;RR#:R0D8_FOoH_OPC05FsRIL_HE80R4-RRI8FMR0FjRR22CRs0MksR8#0_oDFHPO_CFO0s#RH
N
PsLHND#CRk:lRR8#0_oDFHPO_CFO0sL5R_8IH08ERF0IMFRRj2P;
NNsHLRDC8HHP88CMR#:R0D8_FOoH_OPC0RFs5_RNI0H8ERR-4FR8IFM0R2jR;N
PsLHNDsCRCNl_8#[k0RR:#_08DHFoOC_POs0FRL5R_8IH08ERF0IMFRRj2P;
NNsHLRDC0bCl_:LRR8#0_oDFHPO_CFO0sL5R_8IH08ERF0IMFRRj2P;
NNsHLRDCN_bbLRR:#_08DHFoOC_POs0FRL5R_8IH08ERF0IMFRRj2P;
NNsHLRDCs8ClR#:R0D8_FOoH_OPC05FsLH_I8R0E-RR48MFI0jFRRR2;
C
Lo
HM
l#kRR:=50RFE#CsRR=>'Rj'28;
H8PHCRM8:N=R;k
#l25jRR:=N_5NI0H8ERR-4
2;8HHP88CMRR:=8HHP88CM5_RNI0H8ERR-.FR8IFM0R2jRR'&Rj
';N_bbL=R:R''jRR&RL
R;0bCl_:LR=FRM0b5Nb2_LRRR+';4'
l#kRR:=#Rkl+CR0lLb_;H
8PCH8Mj852=R:R0MFR#5RkLl5_8IH0RE22V;
FHsRRRHMjFR0RN5R_8IH0-ERR2.RRFDFbH
SVRR5#5klLH_I820ER'=R42'RRC0EMS
S0bCl_:LR=jR''RR&LS;
CCD#
0SSC_lbL=R:R0MF5bNb_RL2R'+R4
';S8CMR;HV
kS#l=R:Rl#k5IL_HE80R4-RRI8FMR0FjRR2&jR''S;
#5klj:2R=HR8PCH8MR85NH_I8R0E-RR42S;
8HHP88CMRR:=8HHP88CM5_RNI0H8ERR-.FR8IFM0R2jRR'&Rj
';Sl#kRR:=#Rkl+CR0lLb_;8
SH8PHC5M8j:2R=FRM0RR5#5klLH_I820ER
2;CRM8DbFF;V
HR#5RkLl5_8IH0RE2=4R''RR20MEC
CSsl8_N[0k#RR:=#Rkl+RR5'Rj'&RRL2C;
D
#CSlsC_[N8kR#0:#=Rk
l;CRM8H
V;s8ClRR:=s_ClNk8[#R05LH_I8R0E-RR48MFI0jFRR
2;skC0s5MRRP8HHM8C8RR&s8ClRS2;
M
C8HR8P
;
LHCoM-

-kRm00bkR#N#HloMC
M0
FbsO#C#RL5RRL2
CMoH
VSHRL5RRj=R2ER0CSM
SP8HH_8CLj$_RR<=';4'
DSC#SC
SP8HH_8CLj$_RR<=';j'
MSC8VRH;M
C8sRbF#OC#R;RR-

-MRQ0MCsN#DRHNoMD#RN#MHol0CM
s
bF#OC#RR5N
R2LHCoMH
SVRR50lO_FR8C=RR42ER0CSM
SRHV55RNNH_I8R0E-2R4R'=R42'RRC0EMS
SSsbNNRl4<M=RFN052RR+';4'
CSSD
#CSbSSNlsN4=R<R
N;SMSC8VRH;C
SD
#CSNSbs4NlRR<=NS;
CRM8H
V;CRM8bOsFC;##
s
bF#OC#LR52C
Lo
HMSRHV5OR0_8lFCRR=4RR20MEC
HSSVRR5L_5LI0H8ERR-4RR2=4R''RR20MEC
SSSbNNsl<.R=FRM025LR4+R;S
SCCD#
SSSbNNsl<.R=;RL
CSSMH8RVS;
CCD#
bSSNlsN.=R<R
L;S8CMR;HV
8CMRFbsO#C#;


bOsFCR##5NRbs4Nl,NRbs.NlRP2
NNsHLRDCJ0kF_8lFDRR:#_08DHFoOC_POs0FR55RNH_I8R0E+_RLI0H8E-2RR84RF0IMFRRj2
;RLHCoMSS
J0kF_8lFD=R:RP8H5NRbs4Nl,NRbs.NlR
2;SFJk0=R<RFJk0F_l8RD55IN_HE80RL+R_8IH0RE2-84RF0IMF_RLI0H8E;R2
FSl8<DR=kRJFl0_F58DRIL_HE80R4-RRI8FMR0Fj;R2
8CMRFbsO#C#;J

kHF0C_M0.<#R=FRM0k5JFR02+4R''
;

FbsO#C#RJ5Rk,F0RFJk0MHC0#_.,,RNR2LR
oLCHSM
H5VRR55NNH_I8R0E-RR42FRGs5RLLH_I8R0E-RR42=2RR''4R02RE
CMSCS0l<bR=kRJFC0HM.0_#
;RS#CDCS
S0bClRR<=J0kF;SR
CRM8H
V;CRM8bOsFC;##
-

-kRm00bkR#N#HloMC
M0
FbsO#C#RN5RRL,R,FRl82DRSN
PsLHND0CRC4lbR#:R0D8_FOoH_OPC0RFs5_RLI0H8ERR-4FR8IFM0R2jR:5=RREF0CRs#='>R42'R;N
PsLHND0CRC.lbR#:R0D8_FOoH_OPC0RFs5_RNI0H8ERR-4FR8IFM0R2jR;N
PsLHND0CRC.lb_:jRR8#0_oDFHPO_CFO0sRR5NH_I8R0E-RR.8MFI0jFRR=2:RF5R0sEC#>R=R''jR
2;PHNsNCLDRl0Cb:dRR8#0_oDFHPO_CFO0sRR54FR8IFM0R2jR;C
LoRHM
CS0lRbd:N=R5IN_HE80R4-R2RR&L_5LI0H8ERR-4R2;
CS0lRb.:'=R4&'RRl0Cbj._;H
SVRR5s_CllCF8R4=RR02RE
CMSVSHRL5RRj=RR02RE
CMSsSSCHlNMs8CRR<=NL5R_8IH0-ERR84RF0IMFRRj2S;
S#CDH5VRR_0OlCF8R4=RR8NMR=LRRl0CbN4RMN8RR0=RC.lbR02RESCM
SSS-s-RCHlNMs8CRR<=0bCl4S;
SRSRRlsCN8HMC<sR=RR5FC0Es=#R>jR''
2;SDSC#RHV5OR0_8lFCRR=4MRN8RR5lDF8RR/=jRR2NRM8N_5NI0H8ERR-4RR2=4R''RR20MEC
SSSsNClHCM8s=R<R0MF58lFD+2RR''4;S
SCCD#
SSSsNClHCM8s=R<R8lFDS;
S8CMR;HVSSR
CHD#VRR50lO_FR8C=RR42ER0CSM
SVSHRL5RRj=RR02RE
CMSSSSsNClHCM8s=R<RRN5LH_I8R0E-RR48MFI0jFRR
2;SCSSDV#HRL5RR0=RC4lbR8NMR=NRRl0Cb2.RRC0EMS
SS-S-RlsCN8HMC<sR=CR0l;b4
SSSSRRRsNClHCM8s=R<RF5R0sEC#>R=R''jR
2;SCSSD
#CSSSSOCN#R05RCdlbRH2R#SR
SSSSIMECRj"j">R=
SSSSCSslMNH8RCs<l=RF;8DSSR
SSSS
SSSSESIC"MRjR4"=S>
SSSSH5VRR8lFD=R/R2jRRC0EMS
SSSSSsNClHCM8s=R<R+LRR8lFDS;
SSSSCCD#
SSSSsSSCHlNMs8CRR<=lDF8;S
SSCSSMH8RVS;
S
SSSSSSSCIEM4R"j="R>S
SSHSSVRR5lDF8RR/=jRR20MECS
RRSSSSSCSslMNH8RCs<L=RRl-RF;8D
SSSSDSC#SC
SSSSSlsCN8HMC<sR=FRl8
D;SSSSS8CMR;HV
SSSSSS
SSSSIMECR4"4">R=
SSSSVSHRl5RFR8D/j=RR02RE
CMSSSSSCSslMNH8RCs<M=RFl05F28DR'+R4
';SSSSS#CDCS
SSSSSsNClHCM8s=R<R8lFDS;
SSSSCRM8H
V;SSSSSS
SSISSERCMFC0Es=#R>S
SSMSSk;DD
SSSS8CMR#ONCS;
SMSC8VRH;S
SCCD#
SSSH5VRR=LRR2jRRC0EMS
SSCSslMNH8RCs<N=R5_RLI0H8ERR-4FR8IFM0R2jR;S
SS#CDCS
SSCSslMNH8RCs<l=RF;8D
SSSCRM8H
V;SMSC8VRH;

SCRM8bOsFC;##
-
-R0mkbRk0NH##oCMlM
0
bOsFCR##5RRN,,RLRl0CbJ,RkRF02PR
NNsHLRDC0bCl4RR:#_08DHFoOC_POs0FRL5R_8IH0-ERR84RF0IMFRRj2R:=50RFE#CsRR=>'R4'2P;
NNsHLRDC0bCl.RR:#_08DHFoOC_POs0FRN5R_8IH0-ERR84RF0IMFRRj2P;
NNsHLRDC0bCl.R_j:0R#8F_Do_HOP0COF5sRRIN_HE80R.-RRI8FMR0FjRR2:5=RREF0CRs#='>Rj2'R;N
PsLHND0CRCdlbR#:R0D8_FOoH_OPC0RFs5_RNI0H8ERR-4FR8IFM0R2jR;N
PsLHND0CRCdlb_:4RR8#0_oDFHPO_CFO0sRR5NH_I8R0E-RR.8MFI0jFRR:2R=RR5FC0Es=#R>4R'';R2
sPNHDNLCCR0lRbc:0R#8F_Do_HOP0COF5sRRIN_HE80R4-RRI8FMR0Fj:R2=RR5FC0Es=#R>4R'';R2
C
LoRHM
CS0lRb.:'=R4&'RRl0Cbj._;0
SCdlbRR:='Rj'&CR0l_bd4S;
H5VRR/LR=RRj2ER0CSM
S#ONCRR50lO_FR8C2#RH
SSSIMECR=4R>S
SSRHV5RRL=CR0lRb4NRM8NRR=0bCl.RR20MEC
SSSSR--J0kFH0CMRR<=0bCld-;R-HaE#CR)#0kD#MRHR#lHlON0ES
SSRSRRFJk0MHC0=R<Rl0CbR.;
SSSCCD#
SSSSFJk0MHC0=R<Rl0CbS;
SMSC8VRH;S
SSS
SSCIEMRRj=S>
SkSJFC0HM<0R=kRJF
0;S
SSSISSERCMFC0Es=#R>S
SSDMkDS;
SSS
S8CMR#ONCS;
CCD#
OSSNR#C5OR0_8lFCRR2HS#
SESIC4MRR
=>SHSSVRR5N_5NI0H8ERR-4RR2=4R''RR20MEC
SSSSFJk0MHC0=R<Rl0Cb
.;SCSSD
#CSSSSJ0kFH0CMRR<=0bCld
;RSCSSMH8RVR;S
SSS
SSSIMECR=jR>S
SSFJk0MHC0=R<Rl0CbRc;
SSS
SSSIMECREF0CRs#=S>
SkSMD
D;SMSC8NRO#
C;S8CMR;HVSM
C8sRbF#OC#
;
CRM8s;0D
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HON0sHED3NDk;
#HCRC3CC#_08DHFoOM_k#MHoCN83D
D;
0CMHR0$1e7QR
H#RRRRoCCMs5HO
RSRRHRI8R0ERH:RMo0CC:sR=(R4;R
SRsRRI0H8E:RRR0HMCsoCRR:=4
(;SRRRRHNI8R0E:MRH0CCos=R:R
g;SRRRRHLI8R0E:MRH0CCos=R:R;U2
RRRRsbF0S5
R:SqRRHM#_08DHFoOC_POs0F5HNI8R0E-84RF0IMF2Rj;S
SAH:RM0R#8F_Do_HOP0COFLs5I0H8E4R-RI8FMR0Fj
2;SQS7e Q7RF:Rk#0R0D8_FOoH_OPC05FsI0H8E4R-RI8FMR0Fj
2;S S)vhqQ7RS:FRk0#_08DHFoOC_POs0F5HsI8-0E4FR8IFM0R2j2;M
C87R1Q
e;
s
NO0EHCkO0sOCRC_DDDCCPDVRFRQ17e#RH
O
SFFlbM0CMR_7W8
HPSMoCCOsH5S
SNH_I8S0ERm:u1QQae
 ;S_SLI0H8E:SRuQm1a Qe;S
S0lO_FS8CRq:haqz)p
R;SCSslF_l8:CRhzqa)
qpS;S2
FSbs
05SRSNS:SSRRHM#_08DHFoOC_POs0F5IN_HE80-84RF0IMF2Rj;S
SLSRSSH:RM0R#8F_Do_HOP0COFLs5_8IH04E-RI8FMR0Fj
2;SkSJFC0HM:0SR0FkR8#0_oDFHPO_CFO0s_5NI0H8ER-48MFI0jFR2S;
SlsCN8HMC:sSR0FkR8#0_oDFHPO_CFO0s_5LI0H8ER-48MFI0jFR2S;
SP8HH_8CLj$_SF:Rk#0R0D8_FOoH
2SS;C
SMO8RFFlbM0CM;L

CMoH
H
SVC_oMNCs0bC_D:k#RRHV5HNI8R0E>L=RI0H8Eo2RCsMCN
0CS#SSHNoMD_RJNRkGR#:R0D8_FOoH_OPC05FsN8IH0-ER4FR8IFM0R;j2RSR
SHS#oDMNRNs_kRGR:0R#8F_Do_HOP0COFLs5I0H8E4R-RI8FMR0FjR2;RL
SCMoH
lSSk4D0:7RRWH_8PS
SSMoCCOsHRblNRS5
SNSS_8IH0=ER>IRNHE80,S
SS_SLI0H8E>R=RHLI8,0E
SSSS_0OlCF8RR=>4S,
SsSSCll_FR8C=4>R
SSS2S
SSsbF0NRlb
R5SSSSN>R=R
q,SSSSL>R=R
A,SSSSJ0kFH0CMRR=>Jk_NGS,
SsSSCHlNMs8CRR=>sk_NGS
SS
2;S

SSSRSHoV_CsMCN_0C4H:RVsR5I0H8ERR>L8IH0RE2oCCMsCN0
SSSSv) q7QhRR<=15Xask_NGs,RI0H8E
2;SCSSMo8RCsMCNR0CHoV_CsMCN_0C4S;

SSRS_HVoCCMsCN0_R.:H5VRs8IH0<ER=IRLHE802CRoMNCs0SC
S)SS Qvqh<7R=_RsN5kGs8IH04E-RI8FMR0Fj
2;SCSSMo8RCsMCNR0CHoV_CsMCN_0C.S;

SSRS_HVoCCMsCN0_Rd:H5VRI0H8ERR>N8IH0RE2oCCMsCN0
SSSSe7QQR7 <1=RXJa5_GNk,HRI8R0E2S;
SMSC8CRoMNCs0HCRVC_oMNCs0dC_;

SSSRSHoV_CsMCN_0CcH:RVIR5HE80RR<=N8IH0RE2oCCMsCN0
SSSSe7QQR7 <J=R_GNk58IH04E-RI8FMR0Fj
2;SCSSMo8RCsMCNR0CHoV_CsMCN_0CcS;
RMRC8CRoMNCs0HCRVC_oMNCs0bC_D;k#
R
SHoV_CsMCN_0ClkND#H:RVNR5I0H8ERR<L8IH0RE2oCCMsCN0
#SSHNoMD_RNCRG0R#:R0D8_FOoH_OPC05FsL8IH0-ER4FR8IFM0R;j2RRRSSS
S#MHoNJDR_GNkRRR:#_08DHFoOC_POs0F5HLI8R0E-84RF0IMF2Rj;
RRSHS#oDMNRNs_kRGR:0R#8F_Do_HOP0COFLs5I0H8E4R-RI8FMR0FjR2;RR
SLHCoMR
SSCN_G<0R=XR1a,5qRHLI820E;S
Sl0kD4R:R78W_HSP
SCSoMHCsONRlb
R5SSSSNH_I8R0E=L>RI0H8ES,
SLSS_8IH0=ER>IRLHE80,S
SSOS0_8lFC>R=R
4,SSSSs_CllCF8RR=>4S
SSS2
SFSbsl0RN5bR
SSSS=NR>_RNC,G0
SSSS=LR>,RA
SSSSFJk0MHC0>R=RNJ_k
G,SSSSsNClHCM8s>R=RNs_kSG
S;S2
SS

SSRS_HVoCCMsCN0_R4:H5VRs8IH0>ERRHLI820ERMoCC0sNCS
SS S)vhqQ7=R<Ra1X5Ns_kRG,s8IH0;E2
SSSCRM8oCCMsCN0R_HVoCCMsCN0_
4;SR
SSVSH_MoCC0sNC:_.RRHV5HsI8R0E<L=RI0H8Eo2RCsMCN
0CSSSS)q vQRh7<s=R_GNk5HsI8-0E4FR8IFM0R;j2
SSSCRM8oCCMsCN0R_HVoCCMsCN0_
.;SR
SSVSH_MoCC0sNC:_dRRHV58IH0>ERRHLI820ERMoCC0sNCS
SSQS7e Q7RR<=15XaJk_NGI,RHE80R
2;SCSSMo8RCsMCNR0CHoV_CsMCN_0CdS;

SSRS_HVoCCMsCN0_Rc:H5VRI0H8E=R<RHLI820ERMoCC0sNCS
SSQS7e Q7RR<=Jk_NGH5I8-0E4FR8IFM0R;j2
SSSCRM8oCCMsCN0R_HVoCCMsCN0_
c;SCRRMo8RCsMCNR0CHoV_CsMCN_0ClkND#C;
MO8RC_DDDCCPD
;

