--
@ER--a#EHRDVHC#RHRHIs0M0CRRHMNCMRGM0C8RC8ep]7RN0E0NRlbV#Rk0MOH#FM
R--FFM0RHLkDM0H#FRVs$R1MHbDVR$3RCaERlMkCOsHRN#0Ms8N8HR#lNkD0MHFR-
-RObN	CNoR8NMRObN	CNo
R--L$F8RRH#NHPNDDNLCMRFRsNRFD$N0L$RN##HRFVslCRHC
C3-
-
---R-------------------------------------------------------------------------
---R-RR0aHDRCRRRRR:zRhvQ )Ba_17sRNHl0ECO0HRObN	CNoRsVFRM#$0#ECH-#
-RRRRRRRRRRRR:RRRP)C33R4U7R5CRO344cRg2gc
R--RRRRRRRRRRRRR-:
-RRRpsHLNRs$R:RRRHaE#NRbOo	NCER#NRDDLOCRFHlbDRC8HFM0RDNRHNLss#$R$FlLDNHOD
D$-R-RRRRRRRRRRRRR:NRMlRC8Q   3-
-RRRRRRRRRRRRR
R:-R-RRP7CCbDFCRs#: RQ 7 RqR1B10$MEHC##FRWsM	HosRtF,kbR)uqR(4jn
3d-R-RRRRRRRRRRRRR:-
-RuRRkFsb#RCRRRR:a#EHRObN	CNoRV8CH#MCRlMkCOsHRb0$CN#RMN8RsEH0lHC0OkRVMHO0F
M#-R-RRRRRRRRRRRRR:FRVs#RkCHRI0#ER$EM0C##HRF0FDR#3aRIFMCklsRHO0C$b#sRNCCR8VCHM8-:
-RRRRRRRRRRRR:RRRRRRRR-->hRz1hQt R7:ssCbCM#C0z#Rht1QhR 7MLklCHsRMCRPOs0FRsVFl-
-RRRRRRRRRRRRRRR:RRRR->-RRt1Qh: 7RbsCsCC#MR0#NQR1t7h RlMkLRCsHPMRCFO0sFRVs-l
-RRRRRRRRRRRR:RRRCaER#LNCDRCCMlC0$R0bHCR#$R0b1CRap7_mBtQ3-
-RRRRRRRRRRRRRRR:aRECD0CVl0F#R0LHRRH#0NsC0RC8N0#RElCRFR#0#MHoHOVHNRM0L3H0
R--RRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ROPC0#FsRCNsRbsCsCC#M80CRRHM0'IF#FROlCbDl0CMRsVFl-3
-RRRRRRRRRRRR:RRRHaE#NRbOo	NCFROMH0NMF#RPDCsFCN88sRNHl0ECO0HRCFbsFN0sF#RM-
-RRRRRRRRRRRRRRR:0REC1hQt N7RMz8Rht1QhR 70C$b#a3REbCRNNO	oNCRDR#FO0FMN#HM
R--RRRRRRRRRRRRRk:R#kCVD$R0bOCRFCMPsF#HMV#Rk0MOH#FM3-
-RRRRRRRRRRRRR
R:-R-RRRRRRRRRRRRR:VRQR$NMRoNskMlC0FR0RVNRk0MOHRFMHN#RRDMkDsRNs,N$RMNRkRDDNNss$#RH
R--RRRRRRRRRRRRRs:RCs0kMRC85OCGCHb0F,M#RRHVN,M$RCNsR0MFCH8RMP8HHN8kD2D$3-
-RRRRRRRRRRRRR
R:-R-RR0hFCRRRRRRR:FRhRO8CDNNs0MHF#sRFRV8CH0MHH#FMRN#EDLDRCMRHO8DkCH8RMF,Rs-
-RRRRRRRRRRRRRRR:CDGOk88CRFVsl0,RERH#b	NON3oCRCaERObN	CNoRO8CDNNs0MHFRO8CDCNs#-
-RRRRRRRRRRRRRRR:0RECVOkM0MHF#ER0NO0RNLMRC#RkCL8R$RRNks#C3ERaCNRbOo	NCFRL8-$
-RRRRRRRRRRRR:RRRN#EDLDRCFROM8#HC8sCRC0ERsVFlRND8HCVMHH0FFMRVER0CCR#l0NMHRO#F-V
-RRRRRRRRRRRR:RRRH0E#NRbOo	NCa3RFRFD8CCPDCFbsl#RNO$RE#FFCFR0RbHlDCClM00RE-C
-RRRRRRRRRRRR:RRRObN	CNoR8LF$MRHRC0ER#lF0VRCVHHOCRM0lMNMCNsRPDNHNCLDRR0F0lEC3-
-RRRRRRRRRRRRR
R:-R-RRRRRRRRRRRRR:CR)P.3R35cRq3bsRR4.46gg2-
-RRRRRRRRRRRRRRR:aRECVOkM0MHF#3R767,R3Rn,7,3(RU73RC8F#FRM0GRCHR#0H)MRC.PR3
c3-R-RRRRRRRRRRRRR:ERakR#,0#ECCkRVMHO0FRM#NRsCOlFlCCM08kRF0FR0RlOFbRD$IEH0
R--RRRRRRRRRRRRRQ:R R  #M0N88Ns3-
-RRRRRRRRRRRRR
R:---R-------------------------------------------------------------------------
--DsHLNRs$Q   ;#
kC RQ 1 3ap7_mBtQ_n44cD3ND
;
b	NONRoCh zv)_QB1Ra7H
#
R-R-=========================================================================
==R-R-RlhkCOsHRsNsN0$R$RbC8HCVMHH0F
M#R-R-=========================================================================
==
0RR$RbCz h)1emp z7_ht1QhR 7HN#Rs$sNRq5haqz)pNRsMRoC<R>2F1VRaz7_pQmtBR;
Rb0$ChRz)m 1p7e _t1QhR 7HN#Rs$sNRq5haqz)pNRsMRoC<R>2F1VRaz7_pQmtB
;
RDRNHRN#zh_z1hQt H7R#hRz)m 1p7e _1zhQ th7R;
RHNDNz#R_t1QhR 7Hz#Rh1) m pe7Q_1t7h ;R

RL#k0C$bR1zhQ th7#RHR#sCFCDP8hRz)m 1p7e _1zhQ th7R;
RL#k0C$bRt1QhR 7Hs#RCD#FPRC8z h)1emp 17_Q th7
;
R-R-=========================================================================
==R-R-RHqs0CEl0RHOmsbCNs0F#R:
R=--=========================================================================
=
R-R-R:Q8R4q3
VRRk0MOHRFM"#NL"pR5:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7-;R-MRHR8LF$R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pX' aht]R-48MFI0jFR2R3
RR--)kC#DR0:)kC0sRM#0RECNFL#DCk0RDPNkFCRVRRN1hQt P7RCFO0s3RX
R
R-Q-R8q:R3R.
RMVkOF0HM-R""qR5)Rt:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1QhR 7RR=>"lk#H#Mk"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7)5qt 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k0):RCs0kM0#REPCRNCDkRRFV0RECksMN$HRlMRk#FsbCNF0HMMRFRRN
RR--RRRRRRRR1hQt P7RCFO0s)Rqt
3
R-R-============================================================================
R
R-Q-R8q:R3Rd
RMVkOF0HM+R""pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"kbD#
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5Xvq5pp' aht]),R'hp t2a]-84RF0IMF2Rj3R
R-)-RCD#k0q:R8R8#0RIFzQh1t7h ROPC0#FsRN0E0NRl$CRLRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8Rdq3)R
RVOkM0MHFR""+5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Rl1HHsDNRR0FqR3dIsECCRR)HN#RRCFMR0LHR)zh p1me_ 7zQh1t7h 
R
R-Q-R8q:R3
dpRkRVMHO0F"MR+p"5R1:Raz7_pQmtB);RRz:Rh1) m pe7h_z1hQt R72skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RHDlHN0sRF3RqdERICRsCp#RHRFNRMLCRHz0Rh1) m pe7h_z1hQt 
7
R-R-R:Q8Rcq3
VRRk0MOHRFM"R+"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>#R"b#Dk"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7q5vX'5ppt haR],) 'ph]ta2R-48MFI0jFR2R3
RR--)kC#DR0:q#88RF0IRt1QhR 7P0COFRs#00ENR$lNRRLCF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:q)3c
VRRk0MOHRFM"5+"pRR:z h)1emp 17_Q th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR1lNHDsFR0Rcq3RCIEs)CRRRH#LRH0jVRFRMNRFMM-C0oNH3PC
R
R-Q-R8q:R3
cpRkRVMHO0F"MR+p"5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Rl1HHsDNRR0FqR3cIsECCRRpHL#RHj0RRRFVNFRMMC-MoHN0P
C3
-RR-8RQ:3Rq6R
RVOkM0MHFR""+R:5pR)zh p1me_ 7zQh1t7h ;:R)Rahqzp)q2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"kbD#
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R3
RR--)kC#DR0:q#88RRNMzQh1t7h ROPC0,FsRRp,IEH0RMNRFMM-C0oNHRPCQ hat, )R
)3
-RR-8RQ:3RqnR
RVOkM0MHFR""+R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"kbD#
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5p)' aht]R-48MFI0jFR2R3
RR--)kC#DR0:q#88RMNRFMM-C0oNHRPCQ hat, )RRp,IEH0RRNMzQh1t7h ROPC0,FsR
)3
-RR-8RQ:3Rq(R
RVOkM0MHFR""+R:5pRaQh )t ;:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"D#bk;#"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k0q:R8R8#NQMRhta  R),pN5l$CRLR#bFHP0HCsRFRoMCNP0HCR2,0NFRRt1Qh
 7R-R-RRRRRRRRROPC0,FsR
)3
-RR-8RQ:3RqUR
RVOkM0MHFR""+R:5pR)zh p1me_ 71hQt R7;)Q:Rhta  R)2skC0szMRh1) m pe7Q_1t7h RR=>"D#bk;#"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7p 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k0q:R8R8#NQR1t7h ROPC0,FsRRp,0NFRMhRQa  t)),R3R

R=--=========================================================================
==
-RR-8RQ:3RqgR
RVOkM0MHFR""-R,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RlkHM#
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5Xvq5pp' aht]),R'hp t2a]-84RF0IMF2Rj3R
R-)-RCD#k01:RksL0N#O0RF0IR1zhQ th7CRPOs0F#ER0Nl0RNL$RCVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RqgR)
RMVkOF0HM-R""R5p:hRz)m 1p7e _1zhQ th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR1lNHDsFR0Rgq3RCIEs)CRRRH#NMRFCHRL0hRz)m 1p7e _1zhQ th7R

RR--QR8:qp3g
VRRk0MOHRFM"5-"pRR:1_a7ztpmQRB;)RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1HHlDRNs0qFR3IgRECCsRHpR#RRNFRMCLRH0z h)1emp z7_ht1Qh
 7
-RR-8RQ:3Rq4Rj
RMVkOF0HM-R""pR5,:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"H#lM"k#;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5Xvq5pp' aht]),R'hp t2a]-84RF0IMF2Rj3R
R-)-RCD#k01:RksL0N#O0R1NRQ th7CRPOs0F,,R)RFVslMRNFC0EsQR1t7h ROPC0,FsR
p,R-R-RRRRRRRRRN0E0NRl$FRb#L#HDL$RCVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3Rq4
j)RkRVMHO0F"MR-p"5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Rl1HHsDNRR0Fqj34RCIEs)CRRRH#LRH0jVRFRMNRFMM-C0oNH3PC
R
R-Q-R8q:R3p4j
VRRk0MOHRFM"5-"pRR:1_a7ztpmQRB;)RR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR1lNHDsFR0R4q3jERICRsC)#RHR0LHRFjRVRRNM-FMMNCo0CHP3R

RR--QR8:q434
VRRk0MOHRFM"R-"5Rp:z h)1emp z7_ht1Qh; 7)h:Rq)azqRp2skC0szMRh1) m pe7h_z1hQt =7R>lR"H#Mk"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 7p 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k01:RksL0N#O0RMNRFMM-C0oNHRPCQ hat, )RR),VlsFRRNMzQh1t7h ROPC0,FsR
p3
-RR-8RQ:3Rq4R.
RMVkOF0HM-R""pR5:qRhaqz)p);R:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7>R=RH"lM"k#;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt )75'hp t-a]4FR8IFM0R3j2
-RR-CR)#0kD:kR1LN0sOR0#NzMRht1QhR 7P0COFRs,)V,RsRFlNFRMMC-MoHN0PQCRhta  R),p
3
R-R-R:Q8R4q3dR
RVOkM0MHFR""-R:5pR)zh p1me_ 71hQt R7;)Q:Rhta  R)2skC0szMRh1) m pe7Q_1t7h RR=>"H#lM"k#;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R3
RR--)kC#DR0:10kLs0NO#MRNRaQh )t ,,R)RFVslRRN1hQt P7RCFO0sp,R3R

RR--QR8:qc34
VRRk0MOHRFM"R-"5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1QhR 7=">R#MlHk;#"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj3R
R-)-RCD#k01:RksL0N#O0R1NRQ th7CRPOs0F,,R)RFVslMRNRaQh )t ,3Rp
R
R-=-==========================================================================
=
R-R-R:Q8R4q36R
RVOkM0MHFR""*R,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">Rl0kD"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 75pp' aht]'+)pt ha4]-2FR8IFM0R3j2
-RR-CR)#0kD:CRussVFl0#RElCRkHD0bODHNF0HMbRFC0sNHRFMF0MRIzFRht1QhR 7P0COF
s#R-R-RRRRRRRRRN0E0NRl$FRb#L#HDL$RCVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3Rq4Rn
RMVkOF0HM*R""pR5,:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"k#lD;0"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 75pp' aht]'+)pt ha4]-2FR8IFM0R
j2R-R-R#)Ck:D0RDvk0DHbHRC#0RIF1hQt P7RCFO0s0#RERN0lRN$b#F#H$LDRRLCFRV
RR--RRRRRRRR8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R4q3(R
RVOkM0MHFR""*R:5pR)zh p1me_ 7zQh1t7h ;:R)Rahqzp)q2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"lM#k"D0;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt 575p 'ph]ta+pp' aht]2-4RI8FMR0Fj
23R-R-R#)Ck:D0RDvk0DHbHRC#NzMRht1QhR 7P0COFRs,pI,RHR0ENFRMMC-MoHN0PRC
RR--RRRRRRRRQ hat, )RR)3)#RHRMOFP0CsC08RFMRNR1zhQ th7CRPOs0FR
FVR-R-RRRRRRRRRZ1Q 'Rppt haL]RCsVFCkRlDb0HDNHO0MHF3R

RR--QR8:qU34
VRRk0MOHRFM"R*"5Rp:hzqa);qpRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RMk#lD;0"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7)55'hp t+a]) 'ph]ta-R428MFI0jFR2R3
RR--)kC#DR0:v0kDHHbDCN#RMhRz1hQt P7RCFO0s),R,HRI0NERRMMF-oMCNP0HCR
R-R-RRRRRRQRRhta  R),pp3RRRH#OPFMCCs08FR0RRNMzQh1t7h ROPC0RFsFRV
RR--RRRRRRRR1 QZRp)' aht]CRLVCFsRDlk0DHbH0ONH3FM
R
R-Q-R8q:R3
4gRkRVMHO0F"MR*5"Rpz:Rh1) m pe7Q_1t7h ;:R)RaQh )t 2CRs0MksR)zh p1me_ 71hQt =7R>MR"#k#lD;0"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 75pp' aht]'+ppt ha4]-2FR8IFM0R
j2R-R-R#)Ck:D0RDvk0DHbHRC#NQR1t7h ROPC0,FsRRp,IEH0RRNMQ hat, )RR)3)#RH
-RR-RRRRRRRRFROMsPC0RC80NFRRt1QhR 7P0COFFsRVQR1Zp R'hp tRa]LFCVsRC
RR--RRRRRRRRl0kDHHbDOHN0F
M3
-RR-8RQ:3Rq.Rj
RMVkOF0HM*R""pR5:hRQa  t));R:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7>R=R#"M#Dlk0
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt 575) 'ph]ta+p)' aht]2-4RI8FMR0FjR2
RR--)kC#DR0:v0kDHHbDCN#RRt1QhR 7P0COFRs,)I,RHR0ENQMRhta  R),pp3RR
H#R-R-RRRRRRRRRMOFP0CsC08RFRRN1hQt P7RCFO0sVRFRZ1Q 'R)pt haL]RCsVFCR
R-R-RRRRRRlRRkHD0bODHNF0HM
3
R-R-============================================================================
-RR-R
R-R-Rh ma:VRQRO#CFRM8Nksol0CMRRH#xFCsRsVFR""/RCFbsFN0sN,RRP#CC0sH$CRDP
CDR-R-RRRRRRRRF VR)))mRRH#Hk##C
83
-RR-8RQ:3Rq.R4
RMVkOF0HM/R""pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"P8H"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:HR7PCH8#MRNR1zhQ th7CRPOs0F,,RpRRL$N0MFERCszQh1t7h ROPC0,FsR
)3
-RR-8RQ:3Rq.R.
RMVkOF0HM/R""pR5,:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"P8H"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#N1MRQ th7CRPOs0F,,RpRRL$N0MFERCs1hQt P7RCFO0s),R3R

RR--QR8:qd3.
VRRk0MOHRFM"R/"5Rp:z h)1emp z7_ht1Qh; 7RR):hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">RMH#8P
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k07:RH8PHCN#RMhRz1hQt P7RCFO0sp,R,$RLRMNRFMM-C0oNHRPCQ hat, )R
)3R-R-RRRRRRRRRRQVhmm_wQ_Aa)152RR>p 'ph]ta,ER0C)MRRRH#0MskOCN08FR0Rpp' aht]
3
R-R-R:Q8R.q3cR
RVOkM0MHFR""/R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"8M#H;P"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#NFRMMC-MoHN0PQCRhta  R),pL,R$MRNR1zhQ th7CRPOs0F,3R)
-RR-RRRRRRRRVRQR_hmmAw_Q5a1p>2RRp)' aht]0,RERCMp#RHRk0sM0ONC08RF'R)pt ha
]3
-RR-8RQ:3Rq.R6
RMVkOF0HM/R""pR5:hRz)m 1p7e _t1Qh; 7RR):Q hat2 )R0sCkRsMz h)1emp 17_Q th7>R=R#"M#P8H"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:7HHP8RC#NQR1t7h ROPC0,FsRRp,LN$RMhRQa  t)),R3R
R-R-RRRRRRQRRVmRh__mwA1Qa5R)2>'Rppt haR],0MECRH)R#sR0kNMO0RC80pFR'hp t3a]
R
R-Q-R8q:R3
.nRkRVMHO0F"MR/5"RpQ:Rhta  R);)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>MR"#H#8P
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RP7HH#8CRRNMQ hat, )RRp,LN$RRt1QhR 7P0COFRs,)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]RC0EMRRpH0#RsOkMN80CRR0F) 'ph]ta3R

R=--=========================================================================
==R-R-
-RR-hRRm:a RRQV#FCOMN8RslokCRM0Hx#RCRsFVRFs"lsC"bRFC0sNFRs,NCR#PHCs0D$RCDPC
-RR-RRRRRRRRRFV m)))#RHR#H#k3C8
R
R-Q-R8q:R3
.(RkRVMHO0F"MRs"ClR,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RMC#sl
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#Fs3R

RR--QR8:qU3.
VRRk0MOHRFM"lsC"pR5,:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"#M#s"Cl;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0s
#3
-RR-8RQ:3Rq.Rg
RMVkOF0HMsR"CRl"5Rp:z h)1emp z7_ht1Qh; 7RR):hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">RMC#sl
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"spRC)lR"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsNRM8)#RHRRN
RR--RRRRRRRRM-FMMNCo0CHPRaQh )t 3R
R-R-RRRRRRQRRVmRh__mwA1Qa5R)2>'Rppt haR],0MECRH)R#sR0kNMO0RC80pFR'hp t3a]
R
R-Q-R8q:R3
djRkRVMHO0F"MRs"ClR:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"sM#C;l"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRH)R#MRNR1zhQ th7CRPOs0FR8NMRHpR#
RNR-R-RRRRRRRRRMMF-oMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]RC0EMRRpH0#RsOkMN80CRR0F) 'ph]ta3R

RR--QR8:q43d
VRRk0MOHRFM"lsC"pR5:hRz)m 1p7e _t1Qh; 7RR):Q hat2 )R0sCkRsMz h)1emp 17_Q th7>R=R#"M#lsC"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"psRCl)I"RECCsRHpR#QR1t7h ROPC0RFsNRM8)#RHRRNMQ hat3 )
-RR-RRRRRRRRVRQR_hmmAw_Q5a1)>2RRpp' aht]0,RERCM)#RHRk0sM0ONC08RF'Rppt ha
]3
-RR-8RQ:3RqdR.
RMVkOF0HMsR"CRl"5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1QhR 7=">RMs##C;l"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:FRBl0bkC"#RpCRsl"R)RCIEs)CRRRH#1hQt P7RCFO0sMRN8RRpHN#RMhRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]RC0EMRRpH0#RsOkMN80CRR0F) 'ph]ta3R

R=--=========================================================================
==R-R-
-RR-hRRm:a RRQV#FCOMN8RslokCRM0Hx#RCRsFVRFs"8lF"bRFC0sNFRs,NCR#PHCs0D$RCDPC
-RR-RRRRRRRRRFV m)))#RHR#H#k3C8
R
R-Q-R8q:R3
ddRkRVMHO0F"MRl"F8R,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RMF#l8
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#Fs3R

RR--QR8:qc3d
VRRk0MOHRFM"8lF"pR5,:R)R)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0s
#3
-RR-8RQ:3RqdR6
RMVkOF0HMlR"FR8"5Rp:z h)1emp z7_ht1Qh; 7RR):hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">RMF#l8
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsNRM8)R
R-R-RRRRRRHRR#RRNM-FMMNCo0CHPRaQh )t 3R
R-R-RRRRRRQRRVmRh__mwA1Qa5R)2>'Rppt haR],0MECRH)R#sR0kNMO0RC80pFR'hp t3a]
R
R-Q-R8q:R3
dnRkRVMHO0F"MRl"F8R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"lM#F;8"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:BbFlk#0CRR"plRF8)I"RECCsRH)R#MRNR1zhQ th7CRPOs0FR8NMRRp
RR--RRRRRRRRHN#RRMMF-oMCNP0HChRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]RC0EMRRpH0#RsOkMN80CRR0F) 'ph]ta3R

RR--QR8:q(3d
VRRk0MOHRFM"8lF"pR5:hRz)m 1p7e _t1Qh; 7RR):Q hat2 )R0sCkRsMz h)1emp 17_Q th7>R=R#"Ml"F8;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsCp#RHR1NRQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RMhRQa  t)R3
RR--RRRRRRRRQhVRmw_m_aAQ125)Rp>R'hp t,a]RC0EMRR)H0#RsOkMN80CRR0Fp 'ph]ta3R

RR--QR8:qU3d
VRRk0MOHRFM"8lF"pR5:hRQa  t));R:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7>R=R#"Ml"F8;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k0B:RFklb0RC#"lpRF)8R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0sR3
RR--RRRRRRRRQhVRmw_m_aAQ125pR)>R'hp t,a]RC0EMRRpH0#RsOkMN80CRR0F) 'ph]ta3R

R=--=========================================================================
==R-R-R:Q8Rdq3gR
RVOkM0MHFRMVH8C_DVF0l#50RqR)t:hRz)m 1p7e _1zhQ th7Y;RR1:Raz7_pQmtBs2RCs0kMhRQa  t)R;
RR--)kC#D#0Rk$L0bRC:Q hat
 )R-R-R#)Ck:D0RMwH80#REDCRClV0FR#0FkOOsMsCOFCRVER0CNRPDRkCFYVRRRHMq3)t
-RR-RRRRRRRRCR)0Mks#ER0CMRH8RCGF0VREFCROsOksOCMCVRHRRH0C#GH0R#,F-sR40RFEICsH3#C
R
R-Q-R8q:R3
cjRkRVMHO0FVMRH_M8D0CVl0F#R)5qtRR:z h)1emp 17_Q th7Y;RR1:Raz7_pQmtBs2RCs0kMhRQa  t)R;
RR--)kC#D#0Rk$L0bRC:Q hat
 )R-R-R#)Ck:D0RMwH80#REDCRClV0FR#0FkOOsMsCOFCRVER0CNRPDRkCFYVRRRHMq3)t
-RR-RRRRRRRRCR)0Mks#ER0CMRH8RCGF0VREFCROsOksOCMCVRHRRH0C#GH0R#,F-sR40RFEICsH3#C
R
R-Q-R8q:R3
c4RkRVMHO0FVMRH_M8sEHo0#lF0qR5):tRR)zh p1me_ 7zQh1t7h ;RRY:aR17p_zmBtQ2CRs0MksRaQh )t ;R
R-)-RCD#k0kR#Lb0$CQ:Rhta  R)
RR--)kC#DR0:w8HM#ER0CCRDVF0l#F0ROsOksOCMCVRFRC0ERDPNkFCRVRRYHqMR)
t3R-R-RRRRRRRRR0)Ck#sMRC0ER8HMCFGRVER0CORFOsksCCMORRHVHC0RG0H##F,Rs4R-REF0CHsI#
C3
-RR-8RQ:3RqcR.
RMVkOF0HMHRVMs8_H0oEl0F#R)5qtRR:z h)1emp 17_Q th7Y;RR1:Raz7_pQmtBs2RCs0kMhRQa  t)R;
RR--)kC#D#0Rk$L0bRC:Q hat
 )R-R-R#)Ck:D0RMwH80#REDCRClV0FR#0FkOOsMsCOFCRVER0CNRPDRkCFYVRRRHMq3)t
-RR-RRRRRRRRCR)0Mks#ER0CMRH8RCGF0VREFCROsOksOCMCVRHRRH0C#GH0R#,F-sR40RFEICsH3#C
R

R=--=========================================================================
==R-R-RlBFbHNs#RFMmsbCNs0F#R
R-=-==========================================================================
=
R-R-R:Q8R4B3
VRRk0MOHRFM"R>"5Rp,)z:Rh1) m pe7h_z1hQt R72skC0sAMRm mpq=hR>kR"o;0"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R.B3
VRRk0MOHRFM"R>"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph qRR=>"0#o"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCpMRN8RR)NRsC1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RdB3
VRRk0MOHRFM"R>"5Rp:hzqa);qpRR):z h)1emp z7_ht1Qh2 7R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RBcR
RVOkM0MHFR"">R:5pRaQh )t ;:R)R)zh p1me_ 71hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#RRNQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R6B3
VRRk0MOHRFM"R>"5Rp:z h)1emp z7_ht1Qh; 7RR):hzqa)2qpR0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RMhRz1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NFRMMC-MoHN0PQCRhta  
)3
-RR-8RQ:3RBnR
RVOkM0MHFR"">R:5pR)zh p1me_ 71hQt R7;)Q:Rhta  R)2skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#RRN1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NhRQa  t)
3
R-R-============================================================================
R
R-Q-R8B:R3R(
RMVkOF0HM<R""pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qRR=>"0kD"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3RU
RMVkOF0HM<R""pR5,:R)R)zh p1me_ 71hQt R72skC0sAMRm mpq=hR>#R"D;0"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpNRM8)sRNCQR1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3Rg
RMVkOF0HM<R""pR5:qRhaqz)p);R:hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRMNRFMM-C0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:Bj34
VRRk0MOHRFM"R<"5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R4B34R
RVOkM0MHFR""<R:5pR)zh p1me_ 7zQh1t7h ;:R)Rahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-Q-R8B:R3
4.RkRVMHO0F"MR<5"Rpz:Rh1) m pe7Q_1t7h ;:R)RaQh )t 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NQR1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RB4Rd
RMVkOF0HM<R"=5"Rp),R:hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp h>R=RD"kC
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpNRM8)sRNChRz1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R4B3cR
RVOkM0MHFR="<"pR5,:R)R)zh p1me_ 71hQt R72skC0sAMRm mpq=hR>#R"D;C"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRR8NMRN)Rs1CRQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B634
VRRk0MOHRFM""<=R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRMNRFMM-C0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:Bn34
VRRk0MOHRFM""<=R:5pRaQh )t ;:R)R)zh p1me_ 71hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NQR1t7h ROPC03Fs
R
R-Q-R8B:R3
4(RkRVMHO0F"MR<R="5Rp:z h)1emp z7_ht1Qh; 7RR):hzqa)2qpR0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-Q-R8B:R3
4URkRVMHO0F"MR<R="5Rp:z h)1emp 17_Q th7);R:hRQa  t)s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR<=)I"RECCsRHpR#RRN1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NQMRhta  
)3
-RR-============================================================================R

RR--QR8:Bg34
VRRk0MOHRFM"">=R,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMApmm Rqh=">Rk"oC;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
.jRkRVMHO0F"MR>R="5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph qRR=>"C#o"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRNpRM)8RRCNsRt1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB.R4
RMVkOF0HM>R"=5"Rph:Rq)azqRp;)z:Rh1) m pe7h_z1hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RRMMF-oMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRht1QhR 7P0COF
s3
-RR-8RQ:3RB.R.
RMVkOF0HM>R"=5"RpQ:Rhta  R);)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R.B3dR
RVOkM0MHFR=">"pR5:hRz)m 1p7e _1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRHpR#MRNR1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMF-oMCNP0HChRQa  t)
3
R-R-R:Q8R.B3cR
RVOkM0MHFR=">"pR5:hRz)m 1p7e _t1Qh; 7RR):Q hat2 )R0sCkRsMApmm ;qh
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#">pR="R)RCIEspCRRRH#NQR1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RB.R6
RMVkOF0HM=R""pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qRR=>""CJ;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRR8NMRN)RszCRht1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB.Rn
RMVkOF0HM=R""pR5,:R)R)zh p1me_ 71hQt R72skC0sAMRm mpq=hR>CR"J
";R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRNpRM)8RRCNsRt1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB.R(
RMVkOF0HM=R""pR5:qRhaqz)p);R:hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRMNRFMM-C0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR1zhQ th7CRPOs0F3R

RR--QR8:BU3.
VRRk0MOHRFM"R="5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMmRAmqp hR;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8R.B3gR
RVOkM0MHFR""=R:5pR)zh p1me_ 7zQh1t7h ;:R)Rahqzp)q2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NzMRht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFMM-C0oNHRPCQ hat3 )
R
R-Q-R8B:R3
djRkRVMHO0F"MR=5"Rpz:Rh1) m pe7Q_1t7h ;:R)RaQh )t 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NQR1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RBdR4
RMVkOF0HM/R"=5"Rp),R:hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp h>R=RF"M0"CJ;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCpMRN8RR)NRsCzQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
d.RkRVMHO0F"MR/R="5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph qRR=>"0MFC;J"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRR8NMRN)Rs1CRQ th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bd3d
VRRk0MOHRFM""/=R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qRR=>"0MFC;J"
-RR-CR)#0kDRL#k0C$b:mRAmqp hR
R-)-RCD#k0B:RFklb0RC#"/pR="R)RCIEspCRRRH#NFRMMC-MoHN0PQCRhta  N)RMR8
RR--RRRRRRRR)#RHRRNMzQh1t7h ROPC03Fs
R
R-Q-R8B:R3
dcRkRVMHO0F"MR/R="5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMmRAmqp h>R=RF"M0"CJ;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#RRN1hQt P7RCFO0s
3
R-R-R:Q8RdB36R
RVOkM0MHFR="/"pR5:hRz)m 1p7e _1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h>R=RF"M0"CJ;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMzQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNM-FMMNCo0CHPRaQh )t 3R

RR--QR8:Bn3d
VRRk0MOHRFM""/=R:5pR)zh p1me_ 71hQt R7;)Q:Rhta  R)2skC0sAMRm mpq=hR>MR"FJ0C"R;
RR--)kC#D#0Rk$L0bRC:Apmm 
qhR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#RRN1hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NQMRhta  
)3
-RR-============================================================================R

RR--QR8:B(3d
VRRk0MOHRFMvQQhvRzv5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7R
R-)-RCD#k0):RCs0kM0#REDCRCC##sVRFRF0IR)zh p1me_ 7zQh1t7h ROPC0#FsRN0E0NRl$CRL
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBdRU
RMVkOF0HMQRvhzQvvpR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7R
R-)-RCD#k0):RCs0kM0#REDCRCC##sVRFRF0IR)zh p1me_ 71hQt P7RCFO0s0#RERN0lRN$LRC
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bg3d
VRRk0MOHRFMvQQhvRzv5:pRRahqzp)q;RR):hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRRMMFMNCo0CHPRaQh )t ,,RpR8NM
-RR-RRRRRRRRMRNR)zh p1me_ 7zQh1t7h ROPC0,FsR
)3
-RR-8RQ:3RBcRj
RMVkOF0HMQRvhzQvvpR5RQ:Rhta  R);)RR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh
 7R-R-R#)Ck:D0R0)Ck#sMRC0ER#DC#RCsFNVRMhRQa  t)p,R,MRN8MRNR)zh p1me_ 71hQt R7
RR--RRRRRRRRP0COFRs,)
3
R-R-R:Q8RcB34R
RVOkM0MHFRhvQQvvzRR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 
-RR-CR)#0kD:CR)0Mks#ER0CCRD#s#CRRFVNzMRh1) m pe7h_z1hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRRMMFMNCo0CHPRaQh )t ,3R)
R
R-Q-R8B:R3
c.RkRVMHO0FvMRQvhQz5vRpRR:z h)1emp 17_Q th7);RRQ:Rhta  R)2skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 
-RR-CR)#0kD:CR)0Mks#ER0CCRD#s#CRRFVNzMRh1) m pe7Q_1t7h ROPC0,FsRRp,N
M8R-R-RRRRRRRRRRNMQ hat, )R
)3
-RR-============================================================================R

RR--QR8:Bd3c
VRRk0MOHRFMvQqXvRzv5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7R
R-)-RCD#k0):RCs0kM0#REoCRs0CNCFsRVIR0FhRz)m 1p7e _1zhQ th7CRPOs0F#ER0Nl0RNL$RCR
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
ccRkRVMHO0FvMRqvXQz5vRp),RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt R7
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsF0VRIzFRh1) m pe7Q_1t7h ROPC0#FsRN0E0NRl$CRL
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBcR6
RMVkOF0HMqRvXzQvvpR5Rh:Rq)azqRp;)RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7R
R-)-RCD#k0):RCs0kM0#REoCRs0CNCFsRVRRNMMFMC0oNHRPCQ hat, )RRp,N
M8R-R-RRRRRRRRRRNMz h)1emp z7_ht1QhR 7P0COFRs,)
3
R-R-R:Q8RcB3nR
RVOkM0MHFRXvqQvvzRR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt R7
RR--)kC#DR0:)kC0sRM#0RECoNsC0RCsFNVRMhRQa  t)p,R,MRN8MRNR)zh p1me_ 71hQt R7
RR--RRRRRRRRP0COFRs,)
3
R-R-R:Q8RcB3(R
RVOkM0MHFRXvqQvvzRR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 
-RR-CR)#0kD:CR)0Mks#ER0CsRoCCN0sVRFRRNMz h)1emp z7_ht1QhR 7P0COFRs,pN,RMR8
RR--RRRRRRRRNFRMMoMCNP0HChRQa  t)),R3R

RR--QR8:BU3c
VRRk0MOHRFMvQqXvRzv5:pRR)zh p1me_ 71hQt R7;)RR:Q hat2 )R0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7R
R-)-RCD#k0):RCs0kM0#REoCRs0CNCFsRVMRNR)zh p1me_ 71hQt P7RCFO0sp,R,MRN8R
R-R-RRRRRRNRRMhRQa  t)),R3R

R=--=========================================================================
==
-RR-8RQ:3RBcRg
RMVkOF0HM?R">5"Rp),RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRR8NMRN)RszCRh1) m pe7h_z1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R6B3jR
RVOkM0MHFR>"?"pR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCpMRN8RR)NRsCz h)1emp 17_Q th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B436
VRRk0MOHRFM""?>RR5p:qRhaqz)p);RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>"R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7h_z1hQt P7RCFO0s
3
R-R-R:Q8R6B3.R
RVOkM0MHFR>"?"pR5RQ:Rhta  R);)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#">pRRR)"IsECCRRpHN#RRaQh )t R8NM
-RR-RRRRRRRRRR)HN#RMhRz)m 1p7e _t1QhR 7P0COF
s3
-RR-8RQ:3RB6Rd
RMVkOF0HM?R">5"RpRR:z h)1emp z7_ht1Qh; 7R:)RRahqzp)q2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#RpRR>)I"RECCsRHpR#MRNR)zh p1me_ 7zQh1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#RRNMMFMC0oNHRPCQ hat3 )
R
R-Q-R8B:R3
6cRkRVMHO0F"MR?R>"5:pRR)zh p1me_ 71hQt R7;)RR:Q hat2 )R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"R)>R"ERICRsCp#RHRRNMz h)1emp 17_Q th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RB6R6
RMVkOF0HM?R"<5"Rp),RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRR8NMRN)RszCRh1) m pe7h_z1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8R6B3nR
RVOkM0MHFR<"?"pR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"R)<R"ERICRsCpMRN8RR)NRsCz h)1emp 17_Q th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B(36
VRRk0MOHRFM""?<RR5p:qRhaqz)p);RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<"R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7h_z1hQt P7RCFO0s
3
R-R-R:Q8R6B3UR
RVOkM0MHFR<"?"pR5RQ:Rhta  R);)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7Q_1t7h ROPC03Fs
R
R-Q-R8B:R3
6gRkRVMHO0F"MR?R<"5:pRR)zh p1me_ 7zQh1t7h ;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pRRR)"IsECCRRpHN#RMhRz)m 1p7e _1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

RR--QR8:Bj3n
VRRk0MOHRFM""?<RR5p:hRz)m 1p7e _t1Qh; 7R:)RRaQh )t 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#RpRR<)I"RECCsRHpR#MRNR)zh p1me_ 71hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NQMRhta  
)3
-RR-============================================================================R

RR--QR8:B43n
VRRk0MOHRFM"=?<"pR5,RR):hRz)m 1p7e _1zhQ th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRR8NMRN)RszCRh1) m pe7h_z1hQt P7RCFO0sb#RFH##L
D$R-R-RRRRRRRRRRFV8VHVCMsC0CRDMEo0#
3
R-R-R:Q8RnB3.R
RVOkM0MHFR<"?=5"Rp),RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpNRM8)sRNChRz)m 1p7e _t1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RBnRd
RMVkOF0HM?R"<R="5:pRRahqzp)q;RR):hRz)m 1p7e _1zhQ th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NFRMMoMCNP0HChRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7h_z1hQt P7RCFO0s
3
R-R-R:Q8RnB3cR
RVOkM0MHFR<"?=5"RpRR:Q hat; )R:)RR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p<)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR)zh p1me_ 71hQt P7RCFO0s
3
R-R-R:Q8RnB36R
RVOkM0MHFR<"?=5"RpRR:z h)1emp z7_ht1Qh; 7R:)RRahqzp)q2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R<RR)"IsECCRRpHN#RMhRz)m 1p7e _1zhQ th7CRPOs0FR8NM
-RR-RRRRRRRRRR)HN#RRMMFMNCo0CHPRaQh )t 3R

RR--QR8:Bn3n
VRRk0MOHRFM"=?<"pR5Rz:Rh1) m pe7Q_1t7h ;RR):hRQa  t)s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"<pR="R)RCIEspCRRRH#NzMRh1) m pe7Q_1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RBnR(
RMVkOF0HM?R">R="5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRNpRM)8RRCNsR)zh p1me_ 7zQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
nURkRVMHO0F"MR?">=R,5pR:)RR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCpMRN8RR)NRsCz h)1emp 17_Q th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:Bg3n
VRRk0MOHRFM"=?>"pR5Rh:Rq)azqRp;)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR)zh p1me_ 7zQh1t7h ROPC03Fs
R
R-Q-R8B:R3
(jRkRVMHO0F"MR?">=RR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R>RR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7Q_1t7h ROPC03Fs
R
R-Q-R8B:R3
(4RkRVMHO0F"MR?">=RR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p>)=R"ERICRsCp#RHRRNMz h)1emp z7_ht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-8RQ:3RB(R.
RMVkOF0HM?R">R="5:pRR)zh p1me_ 71hQt R7;)RR:Q hat2 )R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR>=)I"RECCsRHpR#MRNR)zh p1me_ 71hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NQMRhta  
)3
-RR-============================================================================R

RR--QR8:Bd3(
VRRk0MOHRFM""?=R,5pR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRNpRM)8RRCNsR)zh p1me_ 7zQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
(cRkRVMHO0F"MR?R="5Rp,)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtBR
R-)-RCD#k0B:RFklb0RC#"=pRRR)"IsECCRRpNRM8)sRNChRz)m 1p7e _t1QhR 7P0COFRs#b#F#H$LD
-RR-RRRRRRRRVRFRV8HVCCsMD0RC0MoE
#3
-RR-8RQ:3RB(R6
RMVkOF0HM?R"=5"RpRR:hzqa);qpR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#RpRR=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR)zh p1me_ 7zQh1t7h ROPC03Fs
R
R-Q-R8B:R3
(nRkRVMHO0F"MR?R="5:pRRaQh )t ;RR):hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR)zh p1me_ 71hQt P7RCFO0s
3
R-R-R:Q8R(B3(R
RVOkM0MHFR="?"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:hzqa)2qpR0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"R)=R"ERICRsCp#RHRRNMz h)1emp z7_ht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-8RQ:3RB(RU
RMVkOF0HM?R"=5"RpRR:z h)1emp 17_Q th7);RRQ:Rhta  R)2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p="R)RCIEspCRRRH#NzMRh1) m pe7Q_1t7h ROPC0RFsN
M8R-R-RRRRRRRRRH)R#MRNRaQh )t 3R

R=--=========================================================================
==
-RR-8RQ:3RB(Rg
RMVkOF0HM?R"/R="5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRNpRM)8RRCNsR)zh p1me_ 7zQh1t7h ROPC0#FsR#bF#DHL$R
R-R-RRRRRRFRRVHR8VsVCCRM0DoCM03E#
R
R-Q-R8B:R3
UjRkRVMHO0F"MR?"/=R,5pR:)RR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCpMRN8RR)NRsCz h)1emp 17_Q th7CRPOs0F#FRb#L#HDR$
RR--RRRRRRRRF8VRHCVVs0CMRMDCo#0E3R

RR--QR8:B43U
VRRk0MOHRFM"=?/"pR5Rh:Rq)azqRp;)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#RRNMMFMC0oNHRPCQ hatR )N
M8R-R-RRRRRRRRRH)R#MRNR)zh p1me_ 7zQh1t7h ROPC03Fs
R
R-Q-R8B:R3
U.RkRVMHO0F"MR?"/=RR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ
-RR-CR)#0kD:FRBl0bkC"#Rp=R/RR)"IsECCRRpHN#RMhRQa  t)MRN8R
R-R-RRRRRR)RRRRH#NzMRh1) m pe7Q_1t7h ROPC03Fs
R
R-Q-R8B:R3
UdRkRVMHO0F"MR?"/=RR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB
RR--)kC#DR0:BbFlk#0CRR"p/)=R"ERICRsCp#RHRRNMz h)1emp z7_ht1QhR 7P0COFNsRMR8
RR--RRRRRRRR)#RHRMNRFCMMoHN0PQCRhta  
)3
-RR-8RQ:3RBURc
RMVkOF0HM?R"/R="5:pRR)zh p1me_ 71hQt R7;)RR:Q hat2 )R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt
QBR-R-R#)Ck:D0RlBFbCk0#pR"RR/=)I"RECCsRHpR#MRNR)zh p1me_ 71hQt P7RCFO0sMRN8R
R-R-RRRRRR)RRRRH#NQMRhta  
)3
R
R-=-==========================================================================R=
RR--1VEH0MRN8FR)0CN0RMwkOF0HMR#
R=--=========================================================================
==
-RR-8RQ:3R14R
RVOkM0MHFRQ1]wpa_ Rwa5tq):hRz)m 1p7e _1zhQ th7B;Rmazh:qRhaqz)ps2RCs0kMhRz)m 1p7e _1zhQ th7>R=RD"#D
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RsuCVlFs#RRN#VEH0C-DVF0RMMRNR1zhQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0R0AHR''j3R
R-a-REBCRmazhRVDC0#lF0HRL0N#RsDCRF3#0
R
R-Q-R81:R3R.
RMVkOF0HM]R1Q_wa)]QtaqR5)Rt:z h)1emp z7_ht1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">R#"sD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NER#H-V0sEHo0MRFRRNMzQh1t7h ROPC0RFsBhmzaHR0l3C#
-RR-RRRRRRRRERaCNRPOCN08FRb#HH0FRM#NRsCVDHDCI8RHR0EARH0'3j'
-RR-RRRRRRRRERaCmRBzRhasEHo0#lF0HRL0N#RsDCRF3#0
R
R-Q-R81:R3Rd
RMVkOF0HM]R1Q_wapa wR)5qtz:Rh1) m pe7Q_1t7h ;mRBz:haRahqzp)q2CRs0MksR)zh p1me_ 71hQt =7R>#R"D;D"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slR#NRE0HV-VDC0MRFR1NRQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0R0AHR''j3R
R-R-RRRRRRaRREBCRmazhRVDC0#lF0HRL0R#,CCGObq0R)pt' ,waRCNsR#DF0
3
R-R-R:Q8Rc13
VRRk0MOHRFM1w]QaQ_)tR]a5tq):hRz)m 1p7e _t1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsMz h)1emp 17_Q th7>R=Rs"#N
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NER#H-V0sEHo0MRFR1NRQ th7CRPOs0FRzBmh0aRH#lC3R
R-R-RRRRRRaRREPCRN0ONCb8RF0#HH#FMRCNsRDVHDRC8IEH0RC0ERVDC0#lF0HRL0q,R)pt' 3wa
-RR-RRRRRRRRERaCmRBzRhasEHo0#lF0HRL0N#RsDCRF3#0
R
R-=-==========================================================================
=
R-R-============================================================================
R
R-Q-R81:R3R6
RMVkOF0HMmR)a qa_wp aqR5)Rt:z h)1emp z7_ht1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">Rs"FD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NFRs0CN0_VDC0VRFRRNMzQh1t7h ROPC0RFsBhmzaHR0l3C#
R
R-Q-R81:R3Rn
RMVkOF0HMmR)a qa_t)Q]5aRq:)tR)zh p1me_ 7zQh1t7h ;mRBz:haRahqzp)q2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"ssF"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slRsNRF00NCH_soRE0FNVRMhRz1hQt P7RCFO0smRBzRha0CHl#
3
R-R-R:Q8R(13
VRRk0MOHRFM)qmaap _ Rwa5tq):hRz)m 1p7e _t1Qh; 7RzBmhRa:hzqa)2qpR0sCkRsMz h)1emp 17_Q th7>R=RF"sD
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k0u:RCFsVsRl#NFRDoNHODFRs0CN0-VDC0VRFR1NRQ th7R
R-R-RRRRRRPRRCFO0smRBzRha0CHl#
3
R-R-R:Q8RU13
VRRk0MOHRFM)qmaa) _Qat]R)5qtz:Rh1) m pe7Q_1t7h ;mRBz:haRahqzp)q2CRs0MksR)zh p1me_ 71hQt =7R>sR"F;s"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:uVCsF#slRDNRFOoHNsDRF00NCH-soRE0FNVRRt1Qh
 7R-R-RRRRRRRRROPC0RFsBhmzaHR0l3C#
R
R-=-==========================================================================R=

-RR-============================================================================

RR-R-----------------------------------------------------------------------------
-RR-RRRhCF0:kRwMHO0F1MR3HgR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-R-RR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rg13
VRRk0MOHRFM"D#D"qR5)Rt:z h)1emp z7_ht1Qh; 7RzBmhRa:Q hat2 )R0sCkRsMz h)1emp z7_ht1QhR 7=">R#"DD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_wp a)5qtB,Rmazh2

RR-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413j#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-RRRFRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1j34
VRRk0MOHRFM"D#D"qR5)Rt:z h)1emp 17_Q th7B;Rmazh:hRQa  t)s2RCs0kMhRz)m 1p7e _t1QhR 7=">R#"DD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]wpa_ 5waq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-R-RR0hFCw:Rk0MOHRFM1434RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-RFRRk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1p08R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:1434
VRRk0MOHRFM"D#s"qR5)Rt:z h)1emp z7_ht1Qh; 7RzBmhRa:Q hat2 )R0sCkRsMz h)1emp z7_ht1QhR 7=">R#"sD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_t)Q]qa5)Rt,BhmzaR2

-RR-----------------------------------------------------------------------------R
R-R-RR0hFCw:Rk0MOHRFM1.34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-RFRRk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4.RkRVMHO0F"MR#"sDR)5qtz:Rh1) m pe7Q_1t7h ;mRBz:haRaQh )t 2CRs0MksR)zh p1me_ 71hQt =7R>#R"s;D"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:z h)1emp 17_Q th7]51Q_wa)]Qtah5z1hQt q75),t2RzBmh2a2
RR
R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1d34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413dR
RVOkM0MHFRF"sD5"Rq:)tR)zh p1me_ 7zQh1t7h ;mRBz:haRaQh )t 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>"DsF"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:)qmaap _ 5waq,)tRzBmh
a2RR
R-----------------------------------------------------------------------------R-
RR--QR8:1c34
VRRk0MOHRFM"DsF"qR5)Rt:z h)1emp 17_Q th7B;Rmazh:hRQa  t)s2RCs0kMhRz)m 1p7e _t1QhR 7=">Rs"FD;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0Ra)mq_a pa w5tq),mRBz2ha
RR
R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1634RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-RFRRk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
46RkRVMHO0F"MRs"FsR)5qtz:Rh1) m pe7h_z1hQt R7;BhmzaQ:Rhta  R)2skC0szMRh1) m pe7h_z1hQt =7R>sR"F;s"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7)5qt 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:mR)a qa_t)Q]qa5)Rt,BhmzaR2

-RR-----------------------------------------------------------------------------R
R-R-RR0hFCw:Rk0MOHRFM1n34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-RFRRk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4nRkRVMHO0F"MRs"FsR)5qtz:Rh1) m pe7Q_1t7h ;mRBz:haRaQh )t 2CRs0MksR)zh p1me_ 71hQt =7R>sR"F;s"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:)qmaa) _Qat]5tq),mRBz2ha
RR
R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFM1(34RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R413(R
RVOkM0MHFRD"#N5"RqR)t:hRz)m 1p7e _1zhQ th7B;RmazhRQ:Rhta  R)2skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]wpa_ 5waq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14HUR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4URkRVMHO0F"MR#"DNR)5qtRR:z h)1emp 17_Q th7B;RmazhRQ:Rhta  R)2skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5tq)'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RQ1]wpa_ 5waq,)tRzBmh
a2
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3R14HgR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R81:R3
4gRkRVMHO0F"MR#"sNR)5qtRR:z h)1emp z7_ht1Qh; 7RzBmh:aRRaQh )t 2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt q75)pt' aht]R-48MFI0jFR2R
R-)-RCD#k01:R]aQw_t)Q]qa5)Rt,Bhmza
2
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR.13j#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R1.Rj
RMVkOF0HM#R"sRN"5tq)Rz:Rh1) m pe7Q_1t7h ;mRBzRha:hRQa  t)s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7q')tpt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1w]QaQ_)t5]aq,)tRzBmh
a2

RRR-R-============================================================================
-RR-)RR Z1Q kRwMHO0F
M#R-R-============================================================================
R
R-Q-R8):R3R4
RMVkOF0HM R)1 QZR)5qtz:Rh1) m pe7Q_1t7h ; RhWQ_1ZR :hzqa)2qpR0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7 5hWQ_1Z4 -RI8FMR0FjR2
RR--)kC#DR0:)QC1ZR #0REC1hQt P7RCFO0s)RqtFR0RC0ERC#bOHHVC18RQ3Z 
-RR-RRRRRRRRFRaRCOsNR0CNNRDssoCROPC0,FsRC0ERIMCRCrDVF0l#R09LRH0bHF#0MHF#R
R-R-RRRRRRNRRsVCRHCDD8HRI00ERE#CRHRoMLRH05tq)'wp aR23WMECRk0sM0ONH,Mo
-RR-RRRRRRRRER0CHR#oLMRHH0R#CRs0MNHCN8RDoFMR0IHEER0CHRsolE0FR#0b0Ns3R

RR--QR8:)
3.RkRVMHO0F)MR Z1Q qR5)Rt:z h)1emp z7_ht1Qh; 7RWh _Z1Q h:Rq)azqRp2skC0szMRh1) m pe7h_z1hQt =7R>0R"s"Hl;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt h75 1W_Q-Z 4FR8IFM0R
j2R-R-R#)Ck:D0R1)CQ#Z RC0ERt1QhR 7P0COFqsR)0tRFER0CbR#CVOHHRC81 QZ3R
R-R-RRRRRRaRRFsROCCN0RDNRNCsosCRPOs0F,ER0CCRMIDRrClV0F9#0R0LHR#bFHF0HMR#
RR--RRRRRRRRNRsCVDHDCI8RHR0E'3j'RCWEMsR0kNMO0oHM,ER0CCRDVF0l#L0RH
0#R-R-RRRRRRRRRCNsRF8sb8bC3R

RMVkOF0HM R)1 QZR)5qt1,RQ_Z )R 1:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1QhR 75Z1Q  _)1C'DMEo0-84RF0IMF2Rj
R
RVOkM0MHFR1) QRZ 5tq),QR1Z) _ :1RR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h RQ51Z) _ D1'C0MoER-48MFI0jFR2


R-R-============================================================================
-RR-FRBMsPC#MHFRMwkOF0HMR#
R=--=========================================================================
==
-RR-8RQ:3R74R
RVOkM0MHFR_amQ hatR )5tq):hRz)m 1p7e _1zhQ th7s2RCs0kMqRhaqz)p>R=Rk"LV;H"
-RR-CR)#0kDRL#k0C$b:qRhaqz)pe3RNCDkRMONMRF0LMCRC0oNHRPC#OHMCNRbsCNl0RCsHN#RMR
R-R-RRRRRRRRRRRRRRzRRht1QhR 7P0COF
s3R-R-R#)Ck:D0RMBFP0Cs#ER0ChRz1hQt P7RCFO0sFR0RRNMQ hat3 )
R
R-Q-R87:R3R.
RMVkOF0HMmRa_aQh )t R)5qtz:Rh1) m pe7Q_1t7h 2CRs0MksRaQh )t RR=>"VLk#;H"
-RR-CR)#0kDRL#k0C$b:hRQa  t)R
R-)-RCD#k0B:RFCMPsR0#NQR1t7h ROPC0RFs0NFRMhRQa  t)
3
R-R-R:Q8Rd73
VRRk0MOHRFMazm_ht1QhR 75tq),QR1ZR :hzqa)2qpR0sCkRsMz h)1emp z7_ht1QhR 7=">R0lsH"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 71 QZ-84RF0IMF2Rj
-RR-CR)#0kD:FRBMsPC0N#RRMMF-oMCNP0HChRQa  t)FR0RRNMzQh1t7h ROPC0RFsIEH0
-RR-RRRRRRRRER0CbR#CVOHHRC81 QZ3R

RMVkOF0HMmRa_t1QhR 75tq)RQ:Rhta  R);1 QZRh:Rq)azqRp2skC0szMRh1) m pe7Q_1t7h RR=>"s#0H;l"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 71 QZ-84RF0IMF2Rj
-RR-CR)#0kD:FRBMsPC0N#RMhRQa  t)FR0RzNRh1) m pe7Q_1t7h ROPC0RFsF0VRE#CRbHCOV8HCRZ1Q 
3
RkRVMHO0FaMRmh_z1hQt 57RqR)t:qRhaqz)p1;RQ_Z )R 1:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 71 QZ_1) 'MDCo-0E4FR8IFM0R
j2
VRRk0MOHRFMa1m_Q th7qR5):tRRaQh )t ;QR1Z) _ :1RR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5Z1Q  _)1C'DMEo0-84RF0IMF2Rj


RR-R-============================================================================
-RR-FRpoNHODbRmC0sNF
s#R-R-============================================================================
R
R-Q-R8p:R3R4
RMVkOF0HMMR"FR0"5Rp:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RM"F0;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0a:RCIslHR#CHCMPsF#HMR

RR--QR8:p
3.RkRVMHO0F"MRN"M8R,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RN"M8;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0e:RCFO0shRq7bRFC0sNH
FM
-RR-8RQ:3RpdR
RVOkM0MHFRs"F"pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h RR=>""Fs;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0e:RCFO0s)RmRCFbsHN0F
M
R-R-R:Q8Rcp3
VRRk0MOHRFM"MMN85"Rp),R:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7>R=RN"MM;8"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7#,RNRlCsoNMC#RNRbHMkp0R
-RR-CR)#0kD:CReOs0FRhhq7bRFC0sNH
FM
-RR-8RQ:3Rp6R
RVOkM0MHFRF"Ms5"Rp),R:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7>R=RF"Ms
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h ,NR#lsCRNCMoRRN#HkMb0
RpR-R-R#)Ck:D0ROeC0RFshRm)FsbCNF0HMR

RR--QR8:p
3nRkRVMHO0F"MRG"FsR,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RG"Fs;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7h_z1hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0e:RCFO0smRX)bRFC0sNH
FM
-RR--RR---------------------------------------------------------------------R-
RR--R0hFCRR:aREC8DCON0sNHRFMNRM8HDlbCMlC0HN0FFMRVER0CGR"M"FsRMVkOF0HM#RH
-RR-#RRbHCOVNHODRD$OlFlCCM08MRk0RHDNI0REEHORl0HCER0C]Re7DpRNkMoNRoCERN#LMCC
-RR-FRRVOVHHDND$8RNFCb08#RNRMOF0MNHHRMo#EkORVNRk0MOH3FMRRq0#EkORbNRF0HM,R
R-R-R0RECVDFDFMIHoFROlMlC0l#RNL$RCCRslCFP8DRNFRMoIEH0RH0E#FRM0CHOR0IHE0Fk
-RR-VRRkEs0C"sRFHVVODHN"NRLD0DF0oHMRRFV0#EHR(4jnR3db	NON3oCRRQ0HR#
RR--RC0ER0HMCRM0F0VRERH#CFVVs00RFsRbF8PHCkR#ONERRMVkOF0HMMRFOHCR0CRLOCFl#R
R-R-RNHPNDDNLCMRHRC0ER7e]p0R#NNM8s
83R-R-R-R----------------------------------------------------------------------R
R-Q-R8p:R3R(
RMVkOF0HMGR"M"FsR,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7=">RGsMF"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh, 7Rl#NCNRsMRoCNH#RM0bkRRp
RR--)kC#DR0:e0COFXsRhRm)FsbCNF0HMR

RR--QR8:p
3URkRVMHO0F"MRM"F0R:5pR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h RR=>"0MF"R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7#,RNRlCsoNMC#RNRbHMkp0R
-RR-CR)#0kD:CRasHlI#HCRMsPC#MHF
R
R-Q-R8p:R3Rg
RMVkOF0HMNR"MR8"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>NR"M;8"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh, 7Rl#NCNRsMRoCNH#RM0bkRRp
RR--)kC#DR0:e0COFqsRhF7RbNCs0MHF
R
R-Q-R8p:R3
4jRkRVMHO0F"MRFRs"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>FR"s
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0e:RCFO0s)RmRCFbsHN0F
M
R-R-R:Q8R4p34R
RVOkM0MHFRN"MMR8"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>MR"N"M8;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h ,NR#lsCRNCMoRRN#HkMb0
RpR-R-R#)Ck:D0ROeC0RFsh7qhRCFbsHN0F
M
R-R-R:Q8R4p3.R
RVOkM0MHFRF"Ms5"Rp),R:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7>R=RF"Ms
";R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt R7,#CNlRMsNoNCR#MRHbRk0pR
R-)-RCD#k0e:RCFO0smRh)bRFC0sNH
FM
-RR-8RQ:3Rp4Rd
RMVkOF0HMGR"FRs"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt =7R>GR"F;s"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh, 7Rl#NCNRsMRoCNH#RM0bkRRp
RR--)kC#DR0:e0COFXsRmF)RbNCs0MHF
R
R-R-R---------------------------------------------------------------------
--R-R-RFRh0:CRRCaERO8CDNNs0MHFR8NMRbHlDCClM00NHRFMF0VRE"CRGsMF"kRVMHO0FHMR#R
R-R-R#ObCHOVHN$DDRlOFl0CMCk8RMD0HRRN0IOEHEHR0l0CREeCR]R7pDoNMkCNoR#ENRCLCMR
R-R-RFHVVODHNDN$R80FbCN8R#FROMH0NMoHMRO#kERRNVOkM0MHF30RqRO#kERRNbMFH0R,
RR--RC0ERDVFDHFIMOoRFCllMR0#lRN$LsCRCPlFCN8RDoFMR0IHEER0HM#RFO0HCHRI0kEF0R
R-R-RV0ksERCs"VFVHNOHDL"RNFDD0M0HoVRFRH0E#jR4(dn3RObN	CNo30RQR
H#R-R-RER0CMRH00CMRRFV0#EHRVCVFRs00bFRsHFP8#CRkROENkRVMHO0FFMRMROCHL0RClOFCR#
RR--RNNPHLDNDHCRMER0C]Re7#pR08NMN3s8
-RR--RR---------------------------------------------------------------------R-
RR--QR8:pc34
VRRk0MOHRFM"FGMs5"Rp),R:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7>R=RM"GF;s"
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh, 7Rl#NCNRsMRoCNH#RM0bkRRp
RR--)kC#DR0:e0COFXsRhRm)FsbCNF0HM


R-R-R:Q8R4p36RR
RMVkOF0HMNR"MR8"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FR7qhRCFbsHN0F
M
R-R-R:Q8R4p3nRR
RMVkOF0HMNR"MR8"5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNR7qhRCFbsHN0F
M
R-R-R:Q8R4p3(RR
RMVkOF0HMFR"s5"RpRR:1_a7ztpmQRB;)RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFsmF)RbNCs0MHF
R
R-Q-R8p:R3R4U
VRRk0MOHRFM""FsRR5p:hRz)m 1p7e _1zhQ th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDs)RmRCFbsHN0F
M
R-R-R:Q8R4p3gRR
RMVkOF0HMMR"N"M8RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0sqRhhF7RbNCs0MHF
R
R-Q-R8p:R3R.j
VRRk0MOHRFM"MMN85"RpRR:z h)1emp z7_ht1Qh; 7R:)RR71a_mzpt2QBR0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNsh7qhRCFbsHN0F
M
R-R-R:Q8R.p34RR
RMVkOF0HMMR"FRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FR)hmRCFbsHN0F
M
R-R-R:Q8R.p3.RR
RMVkOF0HMMR"FRs"5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNR)hmRCFbsHN0F
M
R-R-R:Q8R.p3dRR
RMVkOF0HMGR"FRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FR)XmRCFbsHN0F
M
R-R-R:Q8R.p3cRR
RMVkOF0HMGR"FRs"5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 7zQh1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5pp' aht]R-48MFI0jFR2R
R-)-RCD#k0e:RCFO0sO/1NsDNR)XmRCFbsHN0F
M
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR.p36#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3Rp.
6RRkRVMHO0F"MRGsMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7h_z1hQt R72skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFXsRhRm)FsbCNF0HMR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpn3.RRH#MRF0ObFlNL0HDICRHR0EQ   R810R(4jng-4UR(3BlFlC
M0R-R-R0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVFR Q  0R18jR4(4n-gRU(ObFlNL0HH0DH$R3
R----------------------------------------------------------------------------
--R-R-R:Q8R.p3nRR
RMVkOF0HMGR"M"FsRR5p:hRz)m 1p7e _1zhQ th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDshRXmF)RbNCs0MHF
R
R-Q-R8p:R3R.(
VRRk0MOHRFM"8NM"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFqsRhF7RbNCs0MHF
R
R-Q-R8p:R3R.U
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNqsRhF7RbNCs0MHF
R
R-Q-R8p:R3R.g
VRRk0MOHRFM""FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5)pt ha4]-RI8FMR0FjR2
RR--)kC#DR0:1DONNes/CFO0s)RmRCFbsHN0F
M
R-R-R:Q8Rdp3jRR
RMVkOF0HMFR"s5"RpRR:z h)1emp 17_Q th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNsmF)RbNCs0MHF
R
R-Q-R8p:R3Rd4
VRRk0MOHRFM"MMN85"RpRR:1_a7ztpmQRB;)RR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7) 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:OR1NsDN/OeC0RFsh7qhRCFbsHN0F
M
R-R-R:Q8Rdp3.RR
RMVkOF0HMMR"N"M8RR5p:hRz)m 1p7e _t1Qh; 7R:)RR71a_mzpt2QBR0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'5ppt ha4]-RI8FMR0FjR2
RR--)kC#DR0:e0COF1s/ONNDsqRhhF7RbNCs0MHF
R
R-Q-R8p:R3Rdd
VRRk0MOHRFM"sMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFhsRmF)RbNCs0MHF
R
R-Q-R8p:R3Rdc
VRRk0MOHRFM"sMF"pR5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNhsRmF)RbNCs0MHF
R
R-Q-R8p:R3Rd6
VRRk0MOHRFM"sGF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt )75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0RN1OD/Nse0COFXsRmF)RbNCs0MHF
R
R-Q-R8p:R3Rdn
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2CRs0MksR)zh p1me_ 71hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 71hQt p75'hp t-a]4FR8IFM0R
j2R-R-R#)Ck:D0ROeC0/Fs1DONNXsRmF)RbNCs0MHF
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3Rd(HM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:p(3dRR
RVOkM0MHFRM"GFRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h ;R
R-)-RCD#k0kR#Lb0$Cz:Rh1) m pe7Q_1t7h 5p)' aht]R-48MFI0jFR2R
R-)-RCD#k01:RONNDsC/eOs0FRmXh)bRFC0sNH
FM
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpdHUR#FRM0FROl0bNHCLDR0IHE RQ 1 R048Rj-(n4(gU3FRBlMlC0R
R-F-Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFQsR R  1R084nj(-U4g(FROl0bNHDLHH30$
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3RdU
VRRk0MOHRFM"FGMs5"RpRR:z h)1emp 17_Q th7);RR1:Raz7_pQmtBs2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 7p 'ph]ta-84RF0IMF2Rj
-RR-CR)#0kD:CReOs0F/N1ODRNsX)hmRCFbsHN0F
M
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRdp3g#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpdRg
RMVkOF0HMNR"MR8"5:pRR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB3
-RR-CR)#0kD:CR)#0kDRRFVN'M8HRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHjR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cjRkRVMHO0F"MRM8NM"pR5Rz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVNRMMH8'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3
R
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp34#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcR4
RMVkOF0HMFR"s5"RpRR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB
3RR-R-R#)Ck:D0R#)CkRD0FFVRsM'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp.3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3.R
RVOkM0MHFRF"Ms5"RpRR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB
3RR-R-R#)Ck:D0R#)CkRD0FMVRFHs'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3
R
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3d#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcRd
RMVkOF0HMGR"FRs"5:pRR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtBR;
RR--)kC#D#0Rk$L0bRC:1_a7ztpmQRB3
-RR-CR)#0kD:CR)#0kDRRFVG'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHcR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
ccRkRVMHO0F"MRGsMF"pR5Rz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVMRGFHs'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3
R
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp36#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcR6
RMVkOF0HMNR"MR8"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVMRN8M'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpn3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3nR
RVOkM0MHFRN"MMR8"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVNRMMH8'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3
R
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3(#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcR(
RMVkOF0HMFR"s5"RpRR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQ
B;R-R-R#)CkRD0#0kL$:bCR71a_mzpt3QBRR
R-)-RCD#k0):RCD#k0VRFR'FsHRMoNRDDF0VRELCRHR0#F0VREPCRCFO0s
3R
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHUR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
cURkRVMHO0F"MRM"FsRR5p:hRz)m 1p7e _1zhQ th7s2RCs0kMaR17p_zmBtQ;R
R-)-RCD#k0kR#Lb0$C1:Raz7_pQmtB
3RR-R-R#)Ck:D0R#)CkRD0FMVRFHs'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3
R
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3g#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcRg
RMVkOF0HMGR"FRs"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVFRGsM'HoDRNDVRFRC0ER0LH#VRFRC0EROPC03FsRR

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpj36RRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8R6p3jR
RVOkM0MHFRM"GFRs"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzpt;QB
-RR-CR)#0kDRL#k0C$b:aR17p_zmBtQ3RR
RR--)kC#DR0:)kC#DF0RVMRGFHs'MNoRDFDRVER0CHRL0F#RVER0CCRPOs0F3


R-R-============================================================================
-RR-NRv0ROEwOkM0MHF#R
R-=-==========================================================================
=
R-R-R:Q8R4v3
VRRk0MOHRFM1_a7vBqa]pR5,:R)R71a_mzpt2QBR0sCkRsMApmm ;qh
-RR-CR)#0kD:CR0sRl#ObFlN8sCRsbCR71a_tpmQ4B_4RncHCM0M
0
R-R-R:Q8R.v3
VRRk0MOHRFM1_a7vBqa]pR5,:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k00:RC#slRlOFbCNs8CRbsaR17m_pt_QB4c4nR0HMC
M0
-RR-8RQ:3RvdR
RVOkM0MHFR71a_avqB5]Rp),R:hRz)m 1p7e _t1Qh2 7R0sCkRsMApmm ;qh
-RR-CR)#0kD:CR0sRl#ObFlN8sCRsbCR71a_tpmQ4B_4RncHCM0M
0
R-R-R:Q8R6v3
VRRk0MOHRFM1_a7vBqa]pR5,:R)R71a_mzpt_QBea BmR)2skC0sAMRm mpq
h;R-R-R#)Ck:D0Rs0Cl#IHCFROlsbNHM#FRsbCR71a_tpmQ4B_4RncHCM0M
0
R-R-============================================================================
-RR-sRaNDM#NF0HMkRwMHO0F
M#R-R-============================================================================
R
R-Q-R8a:R3R4
RMVkOF0HMmRa_Rj45R1:z h)1emp z7_ht1Qh; 7RqXvua:17m_ptRQB:'=RjR'2skC0szMRh1) m pe7h_z1hQt =7R>LR"k;V"
-RR-CR)#0kD:CRasHlI#RC,'RE'H0#Rs#NMDCN08FR0R''4R8NMR''DRRH#0MsN#0DNCR8
RR--RRRRRRRR0'FRjR'3QNVRRDPNkFCR0sECRN0EMjR''4|''E|''D|''#RHRkVFM
8,R-R-RRRRRRRRRC0ERsNsNH$R#CR#0FR0R05FE#CsRR=>GblN2N,RMN8RRsINMoHMR
H#R-R-RRRRRRRRR#H#k3C8R)1'NCMoRRH#b#sCCCsP8
3
R-R-R:Q8R.a3
VRRk0MOHRFMajm_41R5:hRz)m 1p7e _t1Qh; 7RqXvua:17m_ptRQB:'=RjR'2skC0szMRh1) m pe7Q_1t7h RR=>"VLk"R;
RR--)kC#DR0:alCsICH#,ER''#RHRN0sMN#D0RC80'FR4N'RM'8RDH'R#sR0NDM#N80C
-RR-RRRRRRRRFR0R''j3VRQRPNRNCDkREF0C0sRERNM'|j''|4''|E''RD'HV#RF8kM,R
R-R-RRRRRR0RRENCRs$sNRRH##RC005FRFC0Es=#R>lRGN,b2R8NMRINRNHsMMHoR#R
R-R-RRRRRRHRR#C#k813R'M)NoHCR#sRbCs#CP3C8
R

RR--QR8:a
3dRkRVMHO0FaMRmj_X41R5Rz:Rh1) m pe7h_z1hQt R72skC0szMRh1) m pe7h_z1hQt 
7;R-R-R#)CkRD0#0kL$:bCR)zh p1me_ 7zQh1t7h 5)1'q ht2R
R-)-RCD#k0a:RCIslH,#CR'']RRH#0MsN#0DNC08RF4R''',RpH'R#sR0NDM#N80CRR0F',j'
-RR-RRRRRRRRMRN8NRPD#kCREF0C0sRERNM'|j''|4''|]''Rp'NRsC0MsN#0DNC08RFXR''
3
R-R-R:Q8Rca3
VRRk0MOHRFMaXm_j54R1RR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 71q')h2t 
-RR-CR)#0kD:CRasHlI#RC,'R]'H0#Rs#NMDCN08FR0R''4,pR''#RHRN0sMN#D0RC80'FRj
',R-R-RRRRRRRRR8NMRDPNkRC#FC0EsER0N'MRj''|4''|]''|pN'Rs0CRs#NMDCN08FR0R''X3R

RR--QR8:a
36RkRVMHO0FaMRmj_X45ZR1RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _1zhQ th7'51)tqh R2
RR--)kC#DR0:alCsICH#,]R''#RHRN0sMN#D0RC80'FR4R','Rp'H0#Rs#NMDCN08FR0R''j,R
R-R-RRRRRRNRRMP8RNCDk#0RFERCs0MENR''j|''4|'']|''p|''ZRCNsRN0sMN#D0RC80'FRX
'3
-RR-8RQ:3RanR
RVOkM0MHFR_amXZj4RR51:hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp 17_Q th7'51)tqh R2
RR--)kC#DR0:alCsICH#,]R''#RHRN0sMN#D0RC80'FR4R','Rp'H0#Rs#NMDCN08FR0R''j,R
R-R-RRRRRRNRRMP8RNCDk#0RFERCs0MENR''j|''4|'']|''p|''ZRCNsRN0sMN#D0RC80'FRX
'3
-RR-8RQ:3Ra(R
RVOkM0MHFR_amz4XjRR51:hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7R;
RR--)kC#D#0Rk$L0bRC:z h)1emp z7_ht1Qh5 71q')h2t 
-RR-CR)#0kD:CRasHlI#RC,'R]'H0#Rs#NMDCN08FR0R''4,pR''#RHRN0sMN#D0RC80'FRj
',R-R-RRRRRRRRR8NMRDPNkRC#FC0EsER0N'MRz''|j''|4''|]''|pN'Rs0CRs#NMDCN08FR0R''X3R

RR--QR8:a
3URkRVMHO0FaMRmX_zj54R1RR:z h)1emp 17_Q th7s2RCs0kMhRz)m 1p7e _t1Qh; 7
-RR-CR)#0kDRL#k0C$b:hRz)m 1p7e _t1Qh5 71q')h2t 
-RR-CR)#0kD:CRasHlI#RC,'R]'H0#Rs#NMDCN08FR0R''4,pR''#RHRN0sMN#D0RC80'FRj
',R-R-RRRRRRRRR8NMRDPNkRC#FC0EsER0N'MRz''|j''|4''|]''|pN'Rs0CRs#NMDCN08FR0R''X3R

RR--QR8:a
3gRkRVMHO0FQMR1R_X5:1RR)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph q;R
R-)-RCD#k0kR#Lb0$CA:Rm mpqRh
RR--)kC#DR0:a )zRRHV1FROMH0NMN#RR''z|''X|''Z|''W|''-RDPNkRC,w1qp 0RFEICsH3#C
R
R-Q-R8a:R3
4jRkRVMHO0FQMR1R_X5:1RR)zh p1me_ 71hQt R72skC0sAMRm mpq
h;R-R-R#)CkRD0#0kL$:bCRmAmph q
-RR-CR)#0kD:)RazH RVRR1O0FMN#HMR'NRz''|X''|Z''|W''|-P'RNCDk,qRwpR1 FC0Es#IHC
3
RRRR-=-==========================================================================R=
RR--#H0sMOoRFCMPsF#HMMRN8sRIHR0CFsbCNF0HMR#
R=--=========================================================================
==R-R-RC0ERDVFDHFIMFoRbNCs0MHF#sRNCsRbCV8CH8MC
R
RVOkM0MHFR_0F#H0sM5oRPkNDCRR:z h)1emp z7_ht1Qh2 7R0sCkRsM1Qa)h
t;RkRVMHO0F0MRF0_#soHMRN5PDRkC:hRz)m 1p7e _t1Qh2 7R0sCkRsM1Qa)h
t;
RRRR-------------------------------------------------------------------RRRR
-RR-mRa_)1aQRht5RNMNNDH#NROD8DCRF"0_0L#soHM"#RHRFbsPCH82R
R-----------------------------------------------------------------R--R
R
R-R-RbCGDHHO0RD$8HCVMRC8FsbCNF0HM
#
RDRNHRN#0LF_#H0sMHoR#FR0_s#0HRMor)zh p1me_ 7zQh1t7h R0sCkRsM1Qa)h;t9
NRRD#HNR_0FLs#0HRMoH0#RF0_#soHMRhrz)m 1p7e _t1QhR 7skC0s1MRah)Qt
9;RDRNHRN#0LF_HsMN$0_#soHMRRH#0#F_0MsHozRrh1) m pe7h_z1hQt s7RCs0kMaR1)tQh9R;
RHNDN0#RFH_LM$Ns_s#0HRMoH0#RF0_#soHMRhrz)m 1p7e _t1QhR 7skC0s1MRah)Qt
9;
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:z h)1emp z7_ht1Qh2 7R0sCkRsM1Qa)h
t;RkRVMHO0F0MRF#_F0MsHoPR5NCDkRz:Rh1) m pe7Q_1t7h 2CRs0MksR)1aQ;ht
NRRD#HNR_0FFNO0D0_#soHMRRH#0FF_#H0sMroRz h)1emp z7_ht1QhR 7skC0s1MRah)Qt
9;RDRNHRN#0FF_OD0N_s#0HRMoH0#RF#_F0MsHozRrh1) m pe7Q_1t7h R0sCkRsM1Qa)h;t9
R
RVOkM0MHFR_0FEs#0HRMo5DPNk:CRR)zh p1me_ 7zQh1t7h 2CRs0MksR)1aQ;ht
VRRk0MOHRFM0EF_#H0sM5oRPkNDCRR:z h)1emp 17_Q th7s2RCs0kMaR1)tQh;R
RNNDH#FR0_GEC_s#0HRMoH0#RF#_E0MsHozRrh1) m pe7h_z1hQt s7RCs0kMaR1)tQh9R;
RHNDN0#RFC_EG0_#soHMRRH#0EF_#H0sMroRz h)1emp 17_Q th7CRs0MksR)1aQ9ht;


CRM8h zv)_QB1;a7
H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
ObN	CNoR8LF$zRhvQ )Ba_17#RH
R
R-M-RkRDDsoNMCsRNsRN$O#FM00NM#R

RMOF#M0N0qRhzRR:z h)1emp z7_ht1QhR 758jRF0IMF2R4RR:=5EF0CRs#='>Rj;'2
ORRF0M#NRM0hRq1:hRz)m 1p7e _t1QhR 758jRF0IMF2R4R:RR=FR50sEC#>R=R''j2
;
R-R-RbHlDCClM00NHRFMO0FMs#FD
R
RO#FM00NMR_hmWhq)QRht:mRAmqp h=R:RDVN#RC;RR--8NCVkRD00CFRlRH0IMNsH#Mo
R
R-=-R========================pNFODkR1LFbsolsN#=R==============================
==
VRRk0MOHRFM1hQt h7_zAv_QRa15tq)RQ:Rhta  R)2skC0shMRq)azqHpR#R
RRNRPsLHNDhCRA1QaRh:Rq)azq
p;RRRRPHNsNCLDRRhRR:RRRahqzp)q;R
RLHCoMR
RRVRHRtq)RR>=jER0CRM
RRRRR:hR=)RqtR;
RCRRD
#CRRRRRRRh:-=R5tq)+;42
RRRR8CMR;HV
RRRRQhAa:1R=;R4
RRRRHIEDhCRRj>RRFDFbR
RRRRRhaAQ1=R:RQhAa41+;R
RRRRRh=R:R/hRR
.;RRRRCRM8DbFF;R
RRCRs0MksRQhAa
1;RMRC8kRVMHO0F1MRQ th7z_hvQ_Aa
1;
VRRk0MOHRFMzQh1t7h _vhz_aAQ1qR5):tRRahqzp)q2CRs0MksRahqzp)qR
H#RRRRPHNsNCLDRQhAa:1RRahqzp)q;R
RRNRPsLHNDhCRRRRRRh:Rq)azq
p;RCRLo
HMRRRRh=R:Rtq);R
RRARhQRa1:4=R;R
RRERIHRDChRR>4FRDFRb
RRRRRQhAa:1R=ARhQ+a14R;
RRRRR:hR=RRh/;R.
RRRR8CMRFDFbR;
RsRRCs0kMARhQ;a1
CRRMV8Rk0MOHRFMzQh1t7h _vhz_aAQ1
;
R-R----------------------------------------------------------------------
-
R-R-RH0E#MRH0MCsNVDRk0MOHRFMObFlk#0CRC0ER8N8HF0HMVRFRF0IR)zh p1me_ 7zQh1t7h 
-RR-HRI0HERM0bkR)Bq)RY
RR--*ER0CIR0FsRNoCklMR0#NRsCF0VRE#CRNRlCDoCM0
E
RkRVMHO0FqMR7z7_ht1QhR 75Rp,)RR:z h)1emp z7_ht1Qh; 7R:BRR71a_tpmQ
B2RRRRskC0szMRh1) m pe7h_z1hQt R7
R
H#RRRRO#FM00NMRpp_ Rwa:hRQa  t)RRR:p=R'MDCo-0E4R;
RNRRD#HNRRXpRRRRR:RRR)zh p1me_ 7zQh1t7h 5pp_ Rwa8MFI0jFR2#RHR
p;RRRRNNDH#)RXRRRRRRRR:hRz)m 1p7e _1zhQ th7_5ppa wRI8FMR0FjH2R#;R)
RRRRsPNHDNLC R)1azpRz:Rh1) m pe7h_z1hQt p75_wp aFR8IFM0R;j2
RRRRsPNHDNLCARBQRaRR1:Rap7_mBtQRR:=BR;
RoLCHRM
RVRRFQsRRRHMjFR0Rpp_ RwaDbFF
RRRR)RR p1za25QRR:=BaAQRsGFR5XpQG2RFXsR)25Q;R
RRRRRBaAQRRRRR=R:RA5BQNaRMX8Rp25Q2sRFRA5BQNaRMX8R)25Q2sRFRp5X5RQ2NRM8XQ)52
2;RRRRCRM8DbFF;R
RRCRs0MksR1) z;pa
CRRMV8Rk0MOHRFMq_77zQh1t7h ;R

RR--0#EHR0HMCNsMDkRVMHO0FOMRFklb0RC#0RECNH880MHFRRFV0RIFz h)1emp 17_Q th7R
R-I-RHR0EHkMb0qRB)
)YR-R-R0*RE0CRINFRslokC#M0RCNsRRFV0REC#CNlRMDCo
0E
VRRk0MOHRFMq_771hQt 57Rp),RRz:Rh1) m pe7Q_1t7h ;RRB:aR17m_pt2QB
RRRR0sCkRsMz h)1emp 17_Q th7R
RHR#
RORRF0M#NRM0p _pw:aRRaQh )t R:RR='RpDoCM04E-;R
RRDRNHRN#XRpRRRRRRRR:z h)1emp 17_Q th7_5ppa wRI8FMR0FjH2R#;Rp
RRRRHNDNX#R)RRRRRRRRz:Rh1) m pe7Q_1t7h 5pp_ Rwa8MFI0jFR2#RHR
);RRRRPHNsNCLDR1) zRpa:hRz)m 1p7e _t1Qh5 7p _pw8aRF0IMF2Rj;R
RRNRPsLHNDBCRARQaRRR:1_a7pQmtB=R:R
B;RCRLo
HMRRRRVRFsQMRHR0jRF_Rppa wRFDFbR
RRRRR)z 1pQa52=R:RQBAaFRGspRX5RQ2GRFsXQ)52R;
RRRRRQBAaRRRR:RR=BR5ARQaNRM8XQp52F2RsBR5ARQaNRM8XQ)52F2RsXR5p25QR8NMR5X)Q;22
RRRR8CMRFDFbR;
RsRRCs0kM R)1azp;R
RCRM8VOkM0MHFR7q7_t1Qh; 7
R
R-----------------------------------------------------------------------------R

RR--0#EHR0HMCNsMDsRbF8OCkRsCObFlk#0CR1zhQ th7HR8PHH#FRM
RR--oHHPM0oREJCRkHF0CRM0NRM8sNClHCM8sR3
RFbsOkC8s7CRQmev7hR5zRv,Xh7 m:vRR)zh p1me_ 7zQh1t7h ;R
RRRRRRRRRRRRRRRRRRTRXz,maR X)vhqQRF:Rkz0Rh1) m pe7h_z1hQt R72HR#
RPRRNNsHLRDCau vR:RRR)zh p1me_ 7zQh1t7h 5vhz'MDCoR0E8MFI0jFR2R;
RPRRNNsHLRDCTazmR:RRR)zh p1me_ 7zQh1t7h 5XvqQvvz5vhz'MDCo,0ER X7h'mvDoCM0-E24R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2R;
RNRRD#HNRh7 mRvRR:RRR)zh p1me_ 7zQh1t7h 5 X7h'mvDoCM04E-RI8FMR0FjH2R#7RX vhm;R
RRNRPsLHNDaCRmQuAaRR:Q hat; )
LRRCMoH
RRRRva uRRR:"=Rjh"&z
v;RRRRTazmR:RR=FR50sEC#>R=R''j2R;
RaRRmQuAa=R:R;-4
RRRRsVFRHKRM R7h'mvsoNMCFRDFRb
RRRRRRHV7m hv25KR'=R40'RE
CMRRRRRRRRaAmuQ:aR=;RK
RRRRRRRRHCG0R;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RNRR#s#C0mRauaAQRR>=jCRsb0FsRz"hvQ )Ba_17Q37e7vm:QR7ev,RmR7,F)sR LvR$CRxs
F"RRRRRCR#PHCs0C$RsssF;R

RVRRFKsRRRHMh'zvDoCM05E-aAmuQ4a+2FR8IFM0RDjRF
FbRRRRRVRHRva um5auaAQ+4K+RI8FMR0FK>2R=jR"" &7h5mvaAmuQ8aRF0IMF2RjRC0EMR
RRRRRR Ravau5mQuAa++K4FR8IFM0RRK2:5=Rau v5uamA+QaKR+48MFI0KFR2R2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-j5"" &7h5mvaAmuQ8aRF0IMF2Rj2R;
RRRRRTRRz5maK:2R=4R''R;
RRRRR8CMR;HV
RRRRNRR#s#C0 Ravau5mQuAa++K4=2RR''j
RRRRRRRRbsCFRs0"vhz B)Q_71a3e7Qv:m7R0HMCNsMDsRCsRFsH0MRE8CRH#PHHRFMNFDosEH0lR"
RRRRR#RRCsPCHR0$CFsssR;
RCRRMD8RF;Fb
RRRRzXTmRaRRR:=)Q 1ZT 5z,maRzXTmDa'C0MoE
2;RRRRXv) qRQh:)=R Z1Q  5avRu,Xv) q'QhDoCM0;E2
CRRMb8RsCFO8CksRe7Qv;m7
R
R-----------------OpFN1DRksLbFNosl-#RRH#EVs0/F00NCbRF#------------------------
-
RkRVMHO0FXMR1Rpp5tq)R1:Raz7_pQmtB _eB)am;mRBzRha:qRhaqz)pR2
RsRRCs0kMaR17p_zmBtQ_Be a
m)R#RH
RRRRMOF#M0N0)RqtR_pRQ:Rhta  R)RRRRRRRRRRRRRRRRRRRRRRRRRRR:=q')tDoCM04E-;R
RRDRNHRN#Xtq)RRRRRRR:1_a7ztpmQeB_ mBa))5qtR_p8MFI0jFR2#RHRtq);R
RRNRPsLHND)CR p1zaRR:1_a7ztpmQeB_ mBa))5qtR_p8MFI0jFR2=R:R05FE#CsRR=>'2j';R
RLHCoMR
RRVRHRzBmh<aR=)RqtR_p0MEC
RRRR)RR p1za)5qtR_p8MFI0BFRmazh2=R:R)Xqt)5qt-_pBhmzaFR8IFM0R;j2
RRRR8CMR;HV
RRRR0sCkRsM)z 1p
a;RMRC8kRVMHO0FXMR1;pp
R
RVOkM0MHFR)X1pqR5):tRR71a_mzpt_QBea BmR);BhmzaRR:hzqa)2qp
RRRR0sCkRsM1_a7ztpmQeB_ mBa)R
RHR#
RORRF0M#NRM0q_)tp:RRRaQh )t RRRRRRRRRRRRRRRRRRRRRRRRR:RR=)RqtC'DMEo0-
4;RRRRNNDH#qRX)RtRRRRR:aR17p_zmBtQ_Be a5m)q_)tpFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)q_)tpFR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRHBVRmazhRR<=q_)tpER0CRM
RRRRR1) z5paq_)tpm-BzRha8MFI0jFR2=R:R)Xqt)5qtR_p8MFI0BFRmazh2R;
RCRRMH8RVR;
RsRRCs0kM R)1azp;R
RCRM8VOkM0MHFR)X1p
;
RkRVMHO0FXMR1R)q5tq)R1:Raz7_pQmtB _eB)am;mRBzRha:qRhaqz)pR2
RsRRCs0kMaR17p_zmBtQ_Be a
m)R#RH
RRRRMOF#M0N0)RqtR_pRQ:Rhta  :)R=)RqtC'DMEo0-
4;RRRRNNDH#qRX)RtRRRRR:aR17p_zmBtQ_Be a5m)q_)tpFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)q_)tpFR8IFM0R;j2
RRRRsPNHDNLCBRXmazhRh:Rq)azq:pR=mRBz;ha
LRRCMoH
RRRRRHV5)5qtC'DMEo0RR<=4F2RsXR5BhmzaRR=jR220MECR0sCkRsMq;)t
RRRR#CDCR
RRRRRH5VRXzBmh>aRRtq)_Rp20MECRmXBzRhaRRRRRRRRR=R:Rtq)_
p;RRRRRMRC8VRH;R
RRRRR)z 1pqa5)pt_-mXBzRha8MFI0jFR2RRRRRRRRRRRR=R:R)Xqt)5qtR_p8MFI0XFRBhmza
2;RRRRR R)1azp5tq)_8pRF0IMFqR5)pt_RX-RBhmzaRR+4R22:5=RFC0Es=#R>qRX)qt5)pt_2
2;RRRRCRM8H
V;RRRRskC0s)MR p1zaR;
R8CMRMVkOF0HM1RX)
q;
VRRk0MOHRFMXp)mR)5qtRR:1_a7ztpmQeB_ mBa)B;RmazhRh:Rq)azq
p2RRRRskC0s1MRaz7_pQmtB _eB)am
HRR#R
RRFROMN#0Mq0R)pt_RRR:Q hatR )RRRRRRRRRRRRRRRRRRRRRRRRR=R:Rtq)'MDCo-0E4R;
RNRRD#HNR)XqtRRRR:RRR71a_mzpt_QBea Bmq)5)pt_RI8FMR0FjH2R#)RqtR;
RPRRNNsHLRDC)z 1p:aRR71a_mzpt_QBea Bmq)5)pt_RI8FMR0Fj:2R=qRX)
t;RRRRPHNsNCLDRzBmhRav:hRQa  t)R;
RoLCHRM
RBRRmazhv=R:RzBmhlaRF58Rq_)tpRR+4
2;RRRRHBVRmazhv=R/R0jRE
CMRRRRR R)1azp5tq)_8pRF0IMFmRBzvha2=R:R)Xqt)5qt-_pBhmza8vRF0IMF2Rj;R
RRRRR)z 1pBa5mazhvR-48MFI0jFR2RRR:X=Rq5)tq_)tpFR8IFM0Rtq)_Bp-mazhv2+4;R
RRMRC8VRH;R
RRCRs0MksR1) z;pa
CRRMV8Rk0MOHRFMXp)m;R

RMVkOF0HM)RXm5)RqR)t:aR17p_zmBtQ_Be a;m)RzBmh:aRRahqzp)q2R
RRCRs0MksR71a_mzpt_QBea BmR)
R
H#RRRRO#FM00NMRtq)_RpR:hRQa  t)RRRRRRRRRRRRRRRRRRRRRRRRRRR:q=R)Dt'C0MoE;-4
RRRRHNDNX#RqR)tRRRRR1:Raz7_pQmtB _eB)am5tq)_8pRF0IMF2RjRRH#q;)t
RRRRsPNHDNLC R)1azpR1:Raz7_pQmtB _eB)am5tq)_8pRF0IMF2RjRR:=Xtq);R
RRNRPsLHNDBCRmazhvRR:Q hat; )
LRRCMoH
RRRRzBmhRav:B=RmazhR8lFR)5qtR_p+2R4;R
RRVRHRzBmhRav/j=RRC0EMR
RRRRR)z 1pqa5)pt_-zBmhRav8MFI0jFR2RRRRRRR:X=Rq5)tq_)tpFR8IFM0RzBmh2av;R
RRRRR)z 1pqa5)pt_RI8FMR0Fq_)tpm-Bzvha+R42:X=Rq5)tBhmza4v-RI8FMR0Fj
2;RRRRCRM8H
V;RRRRskC0s)MR p1zaR;
R8CMRMVkOF0HM)RXm
);
-RR----------------pNFODkR1LFbsolsN#RR-)NCD0MHFNFDRb-#--------------------------R

R
--R-R-RMtCCDsNR""=RsVFR)zh p1me_ 7zQh1t7h ROPC0#Fs,NR#lDCRC0MoER
R-R-
RMVkOF0HMhRz1hQt  7_TpzqR,5pR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0s1MRaz7_pQmtB _eB)am5Rp2=aR17p_zmBtQ_Be a5m))
2;RMRC8kRVMHO0FzMRht1Qh_ 7 qTzp
;
R-R-
-RR-CRtMNCsD=R""FRVshRz)m 1p7e _t1QhR 7P0COF,s#Rl#NCCRDMEo0
-RR-R
RVOkM0MHFRt1Qh_ 7 qTzppR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMaR17p_zmBtQ_Be a5m)p=2RR71a_mzpt_QBea Bm))52R;
R8CMRMVkOF0HMQR1t7h _z Tq
p;
-RR-R
R-t-RCsMCN"DR<V"RFzsRh1) m pe7h_z1hQt P7RCFO0sR#,#CNlRMDCo
0ER-R-
VRRk0MOHRFMzQh1t7h _1p 1pR5,RR):hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)25pR1<Raz7_pQmtB _eB)am5;)2
CRRMV8Rk0MOHRFMzQh1t7h _1p 1
;
R-R-
-RR-CRtMNCsD<R""kRVMHO0FVMRFzsRh1) m pe7Q_1t7h ROPC0#Fs,NR#lDCRC0MoER
R-R-
RMVkOF0HMQR1t7h _1p 1pR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMApmm RqhHR#
RPRRNNsHLRDCQ ha)ph_Rz:Rh1) m pe7Q_1t7h 50jRF'RpDoCM04E-2R;
RPRRNNsHLRDCQ ha))h_Rz:Rh1) m pe7Q_1t7h 50jRF'R)DoCM04E-2R;
RoLCHRM
RQRRh)a hR_pR:RR=;Rp
RRRRaQh _)h)RRRRR:=)R;
RQRRh)a h5_pj:2R=FRM0hRQah )_jp52R;
RQRRh)a h5_)j:2R=FRM0hRQah )_j)52R;
RsRRCs0kMaR17p_zmBtQ_Be a5m)Q ha)ph_2RR<1_a7ztpmQeB_ mBa)h5Qah )_;)2
CRRMV8Rk0MOHRFM1hQt p7_ ;11
R
R-R-
RR--tCCMsRND""<=RMVkOF0HMFRVshRz)m 1p7e _1zhQ th7CRPOs0F##,RNRlCDoCM0RE
R
--RkRVMHO0FzMRht1Qh_ 7p1 1__m) qTzppR5,RR):hRz)m 1p7e _1zhQ th7R2
RsRRCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsM1_a7ztpmQeB_ mBa)25pRR<=1_a7ztpmQeB_ mBa)25);R
RCRM8VOkM0MHFR1zhQ th7 _p1m1_)T_ z;qp
R
R-R-
RR--tCCMsRND""<=RMVkOF0HMFRVshRz)m 1p7e _t1QhR 7P0COF,s#Rl#NCCRDMEo0
-RR-R
RVOkM0MHFRt1Qh_ 7p1 1__m) qTzppR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMApmm RqhHR#
R-RR-CRhCN8RD#HNC0#RF#RN#CksR8HMC8GRHOsC0MHF
RRRRsPNHDNLChRQah )_:pRR)zh p1me_ 71hQt j75RR0FpC'DMEo0-;42
RRRRsPNHDNLChRQah )_:)RR)zh p1me_ 71hQt j75RR0F)C'DMEo0-;42
LRRCMoH
RRRRaQh _)hpRRRRRRRRRRRRRRRRRRRRRRRRRRR:p=R;R
RRhRQah )_R)RRRRRRRRRRRRRRRRRRRRRRRRRRR:=)R;
RQRRh)a h5_pjR2RRRRRRRRRRRRRRRRRRRRRR=R:R0MFRaQh _)hp25j;R
RRhRQah )_j)52RRRRRRRRRRRRRRRRRRRRRRRRR:=MRF0Q ha))h_5;j2
RRRR0sCkRsM1_a7ztpmQeB_ mBa)h5Qah )_Rp2<1=Raz7_pQmtB _eB)am5aQh _)h)
2;RMRC8kRVMHO0F1MRQ th7 _p1m1_)T_ z;qp
R
R-=-R======================== FGbs80CRMwkOF0HM=#R=========================S

VOkM0MHFRlMkL_CsFLV_H_0#kHM#o8MC5lMkRM:RNs0kNRD2skC0sMMRNs0kNHDR#S
SPHNsNCLDRb0l,kRMlsLC__FVL#H0RM:RNs0kN
D;SoLCHSM
Sb0lRR:=M;kl
MSSkClLsV_F_0LH#=R:R
4;SESIHRDC0Rlb>RR4DbFF
SSSMLklCFs_VH_L0:#R=kRMlsLC__FVL#H0+
4;S0SSl:bR=lR0b;/.
CSSMD8RF;Fb
sSSCs0kMkRMlsLC__FVL#H0;C
SMM8RkClLsV_F_0LH#M_k#MHoC
8;SMVkOF0HMkRMlsLC__FVL#H0_o#HMRC85lMk:MRH0CCoss2RCs0kMNRM0NksD#RH
PSSNNsHLRDCMLklCFs_VH_L0R#:MkN0s;ND
PSSNNsHLRDC0:lbR0MNkDsN;L
SCMoH
0SSl:bR=kRMlS;
SRHVMRkl<RRj0MEC
RSSRb0lRR:=-k5Ml2+4;S
SCRM8H
V;SkSMlsLC__FVL#H0RR:=4S;
SHIED0CRl>bRRDjRF
FbSRSRMLklCFs_VH_L0:#R=kRMlsLC__FVL#H0+
4;SRSR0Rlb:0=Rl/bRR
.;SMSC8FRDF
b;SCSs0MksRlMkL_CsFLV_H;0#
MSC8kRMlsLC__FVL#H0_o#HM;C8
RRRRMVkOF0HMqR"A51"pz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt H7R#S
SPHNsNCLDR#sCk:D0R)zh p1me_ 71hQt p75'MDCo-0E4FR8IFM0R;j2
RRRRoLCHSM
SRHV5pp5'VDC0=2RR''j2ER0CSM
SCSs#0kDRR:=pS;
S#CDCS
SS#sCkRD0:R=RjRR-pS;
S8CMR;HV
RRRRRRRR0sCkRsMskC#D
0;RRRRC;M8
RRRRMVkOF0HMaR17q_vaRB]5Rp,)1:Raz7_pQmtBs2RCs0kMmRAmqp h#RH
PSSNNsHLRDCskC#D:0RRFLFDMCN;S
SPHNsNCLDR#8NE0MFVMFk8RR:LDFFC;NM
CSLo
HMSCSs#0kDRR:=V#NDCS;
S#8NE0MFVMFk8=R:RDVN#
C;SVSHR0MFRR5p=-R''FRRsRR)=-R''02RE
CMS8SSNM#EFF0VkRM8:0=Rs;kC
SSSskC#D:0R=RRp=;R)
CSSMH8RVS;
S0sCkRsM5#sCkRD0F5sRMRF08EN#MVF0F8kM2
2;S8CM;R
RRkRVMHO0F1MRav7_q]aBR,5pRR):z h)1emp z7_ht1Qh2 7R0sCkRsMApmm RqhHS#
SsPNHDNLCCRs#0kDRL:RFCFDN
M;SNSPsLHNDHCRRH:RMo0CC
s;SNSPsLHNDDCRNs,RNRR:z h)1emp z7_ht1Qh5 7pC'DMEo0R4-RRI8FMR0Fj
2;SNSPsLHNDDCRNRH,sRNH:0R#8F_Do;HO
RRRRoLCHSM
SRDN:p=R;S
Ss:NR=;R)
VSSFHsRRRHMjFR0RDp'C0MoERR-4FRDFSb
SNSDH=R:R5DNH
2;SsSSN:HR=NRs5;H2
SSSHMVRF50RDRNH=-R''sRFRHsNR'=R-R'20MEC
SSSS#sCkRD0:5=RDRNH=NRsH
2;SSSSHMV5Fs0RCD#k002RE
CMSSSSS0sCk5sMw1qp 
2;SSSSCRM8H
V;SCSSD
#CSSSSskC#D:0R=sR0k
C;SCSSMH8RVS;
S8CMRFDFbS;
S0sCk5sMa )z2R;
RCRRM
8;RRRRVOkM0MHFR71a_avqB5]Rp),R:hRz)m 1p7e _t1Qh2 7R0sCkRsMApmm RqhHS#
SsPNHDNLCCRs#0kDRL:RFCFDN
M;SNSPsLHNDHCRRH:RMo0CC
s;SNSPsLHNDDCRNs,RNRR:z h)1emp 17_Q th7'5pDoCM0-ERR84RF0IMF2Rj;S
SPHNsNCLDRHDN,NRsHRR:#_08DHFoOR;
RLRRCMoH
DSSN=R:R
p;SNSsRR:=)S;
SsVFRHHRMRRj0pFR'MDCoR0E-RR4DbFF
SSSDRNH:D=RN25H;S
SSHsNRR:=sHN52S;
SVSHR0MFRN5DHRR='R-'FssRN=HRR''-2ER0CSM
SsSSCD#k0=R:RN5DHRR=s2NH;S
SSVSH50MFR#sCk2D0RC0EMS
SSsSSCs0kMq5wp21 ;S
SSMSC8VRH;S
SS#CDCS
SSCSs#0kDRR:=0Csk;S
SS8CMR;HV
CSSMD8RF;Fb
sSSCs0kM)5az; 2
RRRR8CM;R

RVRRk0MOHRFM1_a7vBqa]pR5,:R)R8#0_FkDo_HOP0COFRs2skC0sAMRm mpqHhR#S
SPHNsNCLDR#sCkRD0:FRLFNDCMS;
SsPNHDNLCRRH:MRH0CCosS;
SsPNHDNLCNRD,NRsR#:R0k8_DHFoOC_POs0F5Dp'C0MoERR-4FR8IFM0R;j2
PSSNNsHLRDCD,NHRHsNR#:R0k8_DHFoOR;
RLRRCMoH
DSSN=R:R
p;SNSsRR:=)S;
SsVFRHHRMRRj0pFR'MDCoR0E-RR4DbFF
SSSDRNH:D=RN25H;S
SSHsNRR:=sHN52S;
SVSHR0MFRN5DHRR='R-'FssRN=HRR''-2ER0CSM
SsSSCD#k0=R:RN5DHRR=s2NH;S
SSVSH50MFR#sCk2D0RC0EMS
SSsSSCs0kMq5wp21 ;S
SSMSC8VRH;S
SS#CDCS
SSCSs#0kDRR:=0Csk;S
SS8CMR;HV
CSSMD8RF;Fb
sSSCs0kM)5az; 2
RRRR8CM;R

RVRRk0MOHRFMsHC#x5CRq:)tR)zh p1me_ 71hQt R7;h_ W1 QZ:qRhaqz)ps2RCs0kMhRz)m 1p7e _t1QhR 7HR#
RRRRRRRRRNRRD#HNR0LH#z:Rh1) m pe7Q_1t7h 5tq)'hp t-a]4FR8IFM0RRj2Hq#R)
t;RRRRRRRRRRRRPHNsNCLDR#sCk:D0R)zh p1me_ 71hQt h75 1W_Q-Z 4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RRRRRRRRRRRRO#FM00NMRoNsp:CMRaQh )t RR:=q')tpt ha
];RRRRLHCoMR
RRRRRRRRRRVRHRs5NoMpCRh=R 1W_Q2Z RC0EMR
RRRRRRRRRRRRRRsRRCs0kMHRL0
#;RRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRR#sCkRD0:5=RFC0Es=#R>)Rqt)5qt 'pw2a2;R
RRRRRRRRRRVRHR 5hWQ_1Z< RRR.20MEC
RRRRRRRRRRRRRRRR0sCkRsMskC#D
0;RRRRRRRRRRRRCRM8H
V;
RRRRRRRRRRRRRHV5Wh _Z1Q RR<.sRFRoNspRCM<2R.RC0EMR
RRRRRRRRRRRRRRsRRCs0kMCRs#0kD;R
RRRRRRRRRRDRC#RHV5oNspRCM< RhWQ_1ZR 20MEC
RRRRRRRRRRRRRRRRCRs#0kD5oNsp-CM.FR8IFM0RRj2:L=RH50#NpsoC.M-RI8FMR0Fj
2;RRRRRRRRRRRRCCD#
RRRRRRRRRRRRRRRRCRs#0kD5Wh _Z1Q R-.8MFI0jFR2=R:R0LH# 5hWQ_1Z. -RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRskC0ssMRCD#k0R;
RCRRM
8;
kSVMHO0F"MR<5"Rpz:Rh1) m pe7h_z1hQt R7;)h:Rq)azqRp2skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_#kMHCoM825);S
SHMVRkHlL0>#RRpp' aht]ER0CSM
SCSs0MksRza) S;
S8CMR;HV
sSSCs0kM<R"",5pR_amzQh1t7h 5R),p 'ph]ta2
2;S8CM;S

VOkM0MHFR""<R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0k#_Mo#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0swMRq p1;S
SCRM8H
V;SCSs0MksR""<5_amzQh1t7h 5Rp,) 'ph]ta2),R2S;
C;M8
V
Sk0MOHRFM"R<"5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0##MHoCp852S;
SRHVMLklHR0#>'R)pt ha0]RE
CMSsSSCs0kMRRp<;Rj
CSSMH8RVS;
S0sCkRsM"5<"a1m_Q th7,5pRp)' aht]R2,)
2;S8CMR""<;S

VOkM0MHFR""<5Rp:z h)1emp 17_Q th7);R:hRQa  t)s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0##MHoC)852S;
SRHVMLklHR0#>'Rppt ha0]RE
CMSsSSCs0kMRRj<;R)
CSSMH8RVS;
S0sCkRsM"5<"pa,RmQ_1t7h 5R),p 'ph]ta2
2;S8CMR""<;R

RRRRRMVkOF0HM<R"=5"Rph:Rq)azqRp;)z:Rh1) m pe7h_z1hQt R72skC0sAMRm mpqHhR#R
RRRRRRRRRPHNsNCLDRlMkL#H0:qRhaqz)pR;
RRRRRoLCHRM
RRRRRRRRRkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;p2
HSSVkRMl0LH#RR>) 'ph]taRC0EMS
SS0sCkRsMw1qp S;
S8CMR;HV
sSSCs0kM<R"=a"5mh_z1hQt p75,'R)pt ha,]2R;)2
RRRRCRRM
8;
RRRRVRRk0MOHRFM""<=R:5pRaQh )t ;:R)R)zh p1me_ 71hQt R72skC0sAMRm mpqHhR#R
RRRRRPHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;p2
HSSVkRMl0LH#RR>) 'ph]taRC0EMS
SS0sCkRsMpRR<jS;
S8CMR;HV
sSSCs0kM<R"=a"5mQ_1t7h 5Rp,) 'ph]ta2),R2S;
CRM8""<=;R

RRRRRMVkOF0HM<R"=5"Rpz:Rh1) m pe7h_z1hQt R7;)h:Rq)azqRp2skC0sAMRm mpqHhR#R
RRRRRPHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#M_k#MHoC)852S;
SRHVMLklHR0#>'Rppt ha0]RE
CMSsSSCs0kM)Raz
 ;SMSC8VRH;S
SskC0s"MR<5="pa,Rmh_z1hQt )75,'Rppt ha2]2;C
SM
8;

RRRRRRRkRVMHO0F"MR<R="5Rp:z h)1emp 17_Q th7);R:hRQa  t)s2RCs0kMmRAmqp h#RH
RRRRPRRNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_o#HM5C8)
2;SVSHRlMkL#H0Rp>R'hp tRa]0MEC
SSSskC0sjMRR)<R;S
SCRM8H
V;SCSs0MksR="<",5pR_am1hQt )75,'Rppt ha2]2;C
SM"8R<;="
R

RRRRRMVkOF0HM>R""pR5:hRz)m 1p7e _1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMw1qp S;
S8CMR;HV
sSSCs0kM>R"",5pR_amzQh1t7h 5R),p 'ph]ta2
2;S8CM;S

VOkM0MHFR"">R:5pRahqzp)q;:R)R)zh p1me_ 7zQh1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0k#_Mo#HM5C8p
2;SVSHRlMkL#H0R)>R'hp tRa]0MEC
SSSskC0saMR);z 
CSSMH8RVS;
S0sCkRsM"5>"azm_ht1Qh5 7p),R'hp t2a],2R);C
SM
8;
kSVMHO0F"MR>5"RpQ:Rhta  R);)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0##_HCoM825p;S
SHMVRkHlL0>#RRp)' aht]ER0CSM
SCSs0MksR>pRR
j;SMSC8VRH;S
SskC0s"MR>a"5mQ_1t7h 5Rp,) 'ph]ta2),R2S;
CRM8";>"
V
Sk0MOHRFM"5>"pz:Rh1) m pe7Q_1t7h ;:R)RaQh )t 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0##_HCoM825);S
SHMVRkHlL0>#RRpp' aht]ER0CSM
SCSs0MksR>jRR
);SMSC8VRH;S
SskC0s"MR>p"5,mRa_t1Qh5 7)p,R'hp t2a]2S;
CRM8";>"
R
RRRRRVOkM0MHFR=">"pR5:hRz)m 1p7e _1zhQ th7);R:qRhaqz)ps2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0#kHM#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMw1qp S;
S8CMR;HV
sSSCs0kM>R"=p"5,mRa_1zhQ th7,5)Rpp' aht];22
MSC8
;
SMVkOF0HM>R"=5"Rph:Rq)azqRp;)z:Rh1) m pe7h_z1hQt R72skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_#kMHCoM825p;S
SHMVRkHlL0>#RRp)' aht]ER0CSM
SCSs0MksRza) S;
S8CMR;HV
sSSCs0kM>R"=a"5mh_z1hQt p75,'R)pt ha,]2R;)2
MSC8
;
SMVkOF0HM>R"=5"RpQ:Rhta  R);)z:Rh1) m pe7Q_1t7h 2CRs0MksRmAmph qR
H#SsPNHDNLCkRMl0LH#h:Rq)azq
p;SoLCHSM
SlMkL#H0RR:=MLklCFs_VH_L0##_HCoM825p;S
SHMVRkHlL0>#RRp)' aht]ER0CSM
SCSs0MksR>pRR
j;SMSC8VRH;S
SskC0s"MR>5="a1m_Q th7,5pRp)' aht]R2,)
2;S8CMR=">"
;
SMVkOF0HM>R"=p"5:hRz)m 1p7e _t1Qh; 7RR):Q hat2 )R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#H_#o8MC5;)2
HSSVkRMl0LH#RR>p 'ph]taRC0EMS
SS0sCkRsMjRR>)S;
S8CMR;HV
sSSCs0kM>R"=p"5,mRa_t1Qh5 7)p,R'hp t2a]2S;
CRM8"">=;


SMVkOF0HM=R"":5pR)zh p1me_ 71hQt R7;)Q:Rhta  R)2skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_o#HM5C8)
2;SVSH5lMkL#H0Rp>R'hp t2a]RC0EMS
SS0sCk5sMw1qp 
2;SDSC#SC
SCSs0MksR""=5Rp,a1m_Q th7,5)Rpp' aht];22
CSSMH8RVS;
CRM8";="
SS
VOkM0MHFR""=5Rp:Q hat; )RR):z h)1emp 17_Q th7s2RCs0kMmRAmqp h#RH
NSPsLHNDMCRkHlL0R#:hzqa);qp
CSLo
HMSkSMl0LH#=R:RlMkL_CsFLV_H_0##MHoCp852S;
S5HVMLklHR0#>'R)pt haR]20MEC
SSSskC0swM5q p12S;
S#CDCS
SS0sCkRsM"5=")a,RmQ_1t7h 5Rp,) 'ph]ta2
2;SMSC8VRH;C
SM"8R=
";
RRRRVRRk0MOHRFM"5="pz:Rh1) m pe7h_z1hQt R7;)h:Rq)azqRp2skC0sAMRm mpqHhR#P
SNNsHLRDCMLklH:0#Rahqzp)q;L
SCMoH
MSSkHlL0:#R=kRMlsLC__FVL#H0_#kMHCoM825);S
SHMV5kHlL0>#RRpp' aht]02RE
CMSsSSCs0kMq5wp21 ;S
SCCD#
SSSskC0s"MR=p"5,mRa_1zhQ th7,5)Rpp' aht];22
CSSMH8RVS;
CRM8";="
SS
VOkM0MHFR""=5Rp:hzqa);qpRR):z h)1emp z7_ht1Qh2 7R0sCkRsMApmm RqhHS#
PHNsNCLDRlMkL#H0:qRhaqz)pS;
LHCoMS
SMLklHR0#:M=RkClLsV_F_0LH#M_k#MHoCp852S;
S5HVMLklHR0#>'R)pt haR]20MEC
SSSskC0swM5q p12S;
S#CDCS
SS0sCkRsM"5=")a,Rmh_z1hQt p75,'R)pt ha2]2;S
SCRM8H
V;S8CMR""=;


SMVkOF0HMlR"FR8"5Rp,)z:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt H7R#P
SNNsHLRDCskC#D:0RR)zh p1me_ 71hQt )75'MDCo-0E4FR8IFM0R;j2
NSPsLHNDsCRCHlNMs8CRz:Rh1) m pe7h_z1hQt )75'MDCo-0E4FR8IFM0R;j2
NSPsLHND0CRlRbD:hRz)m 1p7e _1zhQ th7'5pDoCM04E-RI8FMR0Fj
2;SsPNHDNLClR0b:sRR)zh p1me_ 7zQh1t7h 5D)'C0MoER-48MFI0jFR2S;
PHNsNCLDR8IH0REN:MRH0CCos=R:RDp'C0MoES;
PHNsNCLDR8IH0REL:MRH0CCos=R:RD)'C0MoES;
PHNsNCLDRosHEC0MoA:Rm mpq:hR=qRwp;1 
CSLo
HMSVSHR55pp 'pwRa2=4R''02RE
CMS0SSlRbD:k=RMo#HM5C8-;p2
CSSD
#CS0SSlRbD:k=RMo#HM5C8p
2;SMSC8VRH;S
SH5VR)'5)pa w2RR='24'RC0EMS
SSb0ls=R:R#kMHCoM8)5-2S;
SHSsoME0C:oR=)Raz
 ;SDSC#SC
SlS0b:sR=MRk#MHoC)852S;
S8CMR;HV
HSSVR5)=2RjRC0EMS
SS#sCkRD0:5=RFC0Es=#R>jR''
2;SDSC#RCS
SSS-C-slMNH8
CsSsSSCHlNMs8CRR:="lsC"l50b0D,l2bs;S
SSRHVsEHo0oMCR8NMRpp5'wp a'2=40'RE
CMSRSSRlsCN8HMC:sR=jR""C-slMNH8;Cs
SSSCHD#VHRsoME0CNoRMs8RCHlNMs8C/j=""ER0CSM
SRSRsNClHCM8s=R:RlsCN8HMC0s-l;bs
SSSCHD#V5Rpp 'pw=a2'R4'NRM8sNClHCM8s"/=j0"RE
CMSRSSRlsCN8HMC:sR=lR0bss-CHlNMs8C;S
SSMSC8VRH;S
SS#sCkRD0:1=RQ th7C5slMNH82Cs;S
SCRM8H
V;SCSs0MksR#sCk;D0
MSC8lR"F;8"
R
R-Q-R8q:R3
d)RkRVMHO0F"MR+5"RpRR:z h)1emp z7_ht1Qh; 7R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp z7_ht1Qh
 7R#RH
RRRRsPNHDNLC)RXRz:Rh1) m pe7h_z1hQt p75'MDCo-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRXj)52=R:R
);RRRRskC0s5MRpRR+X;)2
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3
dpRkRVMHO0F"MR+5"RpRR:1_a7ztpmQRB;)RR:z h)1emp z7_ht1Qh2 7
RRRR0sCkRsMz h)1emp z7_ht1Qh
 7R#RH
RRRRsPNHDNLCpRXRz:Rh1) m pe7h_z1hQt )75'MDCo-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRXjp52=R:R
p;RRRRskC0s5MRX+pRR;)2
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3
c)RkRVMHO0F"MR+5"RpRR:z h)1emp 17_Q th7);RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _t1Qh
 7R#RH
RRRRsPNHDNLC)RXRz:Rh1) m pe7Q_1t7h 5Dp'C0MoER-48MFI0jFR2=R:R05FE#CsRR=>'2j';R
RLHCoMR
RR)RX5Rj2:)=R;R
RRCRs0MksRR5p+)RX2R;
R8CMRMVkOF0HM+R""
;
R-R-R:Q8Rcq3pR
RVOkM0MHFR""+RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _t1Qh2 7
RRRR0sCkRsMz h)1emp 17_Q th7R
RHR#
RPRRNNsHLRDCX:pRR)zh p1me_ 71hQt )75'MDCo-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRXjp52=R:R
p;RRRRskC0s5MRX+pRR;)2
CRRMV8Rk0MOHRFM";+"
R
R-Q-R8q:R3
g)RkRVMHO0F"MR-5"RpRR:z h)1emp z7_ht1Qh; 7R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp z7_ht1Qh
 7R#RH
RRRRsPNHDNLC)RXRz:Rh1) m pe7h_z1hQt p75'MDCo-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRXj)52=R:R
);RRRRskC0s5MRpRR-X;)2
CRRMV8Rk0MOHRFM";-"
R
R-Q-R8q:R3
gpRkRVMHO0F"MR-5"RpRR:1_a7ztpmQRB;)RR:z h)1emp z7_ht1Qh2 7
RRRR0sCkRsMz h)1emp z7_ht1Qh
 7R#RH
RRRRsPNHDNLCpRXRz:Rh1) m pe7h_z1hQt )75'MDCo-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLo
HMRRRRXjp52=R:R
p;RRRRskC0s5MRX-pRR;)2
CRRMV8Rk0MOHRFM";-"
R
R-Q-R8q:R3)4j
VRRk0MOHRFM"R-"5:pRR)zh p1me_ 71hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7Q_1t7h 
HRR#R
RRNRPsLHNDXCR)RR:z h)1emp 17_Q th7'5pDoCM04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2R;
RoLCHRM
RXRR)25jRR:=)R;
RsRRCs0kMpR5RX-R)
2;RMRC8kRVMHO0F"MR-
";
-RR-8RQ:3Rq4
jpRkRVMHO0F"MR-5"RpRR:1_a7ztpmQRB;)RR:z h)1emp 17_Q th7R2
RsRRCs0kMhRz)m 1p7e _t1Qh
 7R#RH
RRRRsPNHDNLCpRXRz:Rh1) m pe7Q_1t7h 5D)'C0MoER-48MFI0jFR2=R:R05FE#CsRR=>'2j';R
RLHCoMR
RRpRX5Rj2:p=R;R
RRCRs0MksRp5XR)-R2R;
R8CMRMVkOF0HM-R""
;
R-R-R============================================================================R
R-Q-R8q:R3
dgRkRVMHO0FVMRH_M8D0CVl0F#R)5qtRR:z h)1emp z7_ht1Qh; 7R:YRR71a_mzpt2QB
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RVRRFQsRhX7 RRHMq')tsoNMCFRDFRb
RRRRRRHVq5)tQ h7X?2R=RRY0MEC
RRRRRRRR0sCkRsMQ h7XR;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RsRRCs0kM4R-;R
RCRM8VOkM0MHFRMVH8C_DVF0l#
0;
-RR-8RQ:3RqcRj
RMVkOF0HMHRVMD8_ClV0FR#05tq)Rz:Rh1) m pe7Q_1t7h ;RRY:aR17p_zmBtQ2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRRVRFsQ h7XMRHRtq)'MsNoDCRF
FbRRRRRVRHRtq)57Qh RX2?Y=RRC0EMR
RRRRRRCRs0MksR7Qh 
X;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRRskC0s-MR4R;
R8CMRMVkOF0HMHRVMD8_ClV0F;#0
R
R-Q-R8q:R3
c4RkRVMHO0FVMRH_M8sEHo0#lF0qR5):tRR)zh p1me_ 7zQh1t7h ;RRY:aR17p_zmBtQ2R
RRCRs0MksRaQh )t R
H#RCRLo
HMRRRRVRFsQ h7XMRHRtq)'PsCCCs#_MsNoDCRF
FbRRRRRVRHRtq)57Qh RX2?Y=RRC0EMR
RRRRRRCRs0MksR7Qh 
X;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRRskC0s-MR4R;
R8CMRMVkOF0HMHRVMs8_H0oEl0F#;R

RR--QR8:q.3c
VRRk0MOHRFMV8HM_osHEF0l#50RqR)t:hRz)m 1p7e _t1Qh; 7R:YRR71a_mzpt2QB
RRRR0sCkRsMQ hatR )HR#
RoLCHRM
RVRRFQsRhX7 RRHMq')tsCCPs_#CsoNMCFRDFRb
RRRRRRHVq5)tQ h7X?2R=RRY0MEC
RRRRRRRR0sCkRsMQ h7XR;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RsRRCs0kM4R-;R
RCRM8VOkM0MHFRMVH8H_solE0F;#0
R
R-=-R=========================================================================
==
-RR-8RQ:3RBdR(
RMVkOF0HMQRvhzQvvpR5,RR):hRz)m 1p7e _1zhQ th7s2RCs0kMhRz)m 1p7e _1zhQ th7#RH
RRRRMOF#M0N0QR1Z: RRahqzp)qRR:=vQqXv5zvpC'DMEo0,'R)DoCM0;E2
RRRRsPNHDNLCjRp4:RRR)zh p1me_ 7zQh1t7h 5Z1Q R-48MFI0jFR2R;
RPRRNNsHLRDC)Rj4Rz:Rh1) m pe7h_z1hQt 175Q-Z 4FR8IFM0R;j2
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RERCMskC0shMRq
z;RRRRCRM8H
V;RRRRpRj4:a=Rm4_j51) Q5Z p1,RQ2Z ,XR''
2;RRRRH5VRp5j4p'j4D0CV2RR='2X'RC0EMCRs0MksR4pj;R
RRMRC8VRH;R
RRjR)4=R:R_amj)45 Z1Q ,5)RZ1Q R2,'2X';R
RRVRHRj5)4j5)4C'DVR02=XR''02RERCMskC0s)MRj
4;RRRRCRM8H
V;RRRRHzVRht1Qh_ 7p1 154pj,jR)402RE
CMRRRRRCRs0MksR4pj;R
RRDRC#RC
RRRRR0sCkRsM);j4
RRRR8CMR;HV
CRRMV8Rk0MOHRFMvQQhv;zv
R
R-Q-R8B:R3
dURkRVMHO0FvMRQvhQz5vRp),RRz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt H7R#R
RRFROMN#0M10RQRZ :qRhaqz)p=R:RXvqQvvz5Dp'C0MoE),R'MDCo20E;R
RRNRPsLHNDpCRjR4R:hRz)m 1p7e _t1Qh5 71 QZ-84RF0IMF2Rj;R
RRNRPsLHND)CRjR4R:hRz)m 1p7e _t1Qh5 71 QZ-84RF0IMF2Rj;R
RLHCoMR
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MECR0sCkRsMh;q1
RRRR8CMR;HV
RRRR4pjRR:=ajm_4 5)1 QZ5Rp,1 QZ2',RX;'2
RRRRRHV54pj54pj'VDC0=2RR''X2ER0CsMRCs0kMjRp4R;
RCRRMH8RVR;
R)RRj:4R=mRa_5j4)Q 1Z) 5,QR1Z, 2R''X2R;
RHRRV)R5j)45jD4'C2V0R'=RXR'20MECR0sCkRsM);j4
RRRR8CMR;HV
RRRRRHV1hQt p7_ 511p,j4R4)j2ER0CRM
RRRRR0sCkRsMp;j4
RRRR#CDCR
RRRRRskC0s)MRj
4;RRRRCRM8H
V;RMRC8kRVMHO0FvMRQvhQz
v;
-RR-8RQ:3RBdRg
RMVkOF0HMQRvhzQvvpR5Rh:Rq)azqRp;)RR:z h)1emp z7_ht1Qh2 7
RRRR0sCkRsMz h)1emp z7_ht1QhR 7HR#
RoLCHRM
RsRRCs0kMQRvhzQvvm5a_1zhQ th7,5pRD)'C0MoER2,)
2;RMRC8kRVMHO0FvMRQvhQz
v;
-RR-8RQ:3RBcRj
RMVkOF0HMQRvhzQvvpR5RQ:Rhta  R);)RR:z h)1emp 17_Q th7R2
RsRRCs0kMhRz)m 1p7e _t1QhR 7HR#
RoLCHRM
RsRRCs0kMQRvhzQvvm5a_t1Qh5 7p),R'MDCo20E,2R);R
RCRM8VOkM0MHFRhvQQvvz;R

RR--QR8:B43c
VRRk0MOHRFMvQQhvRzv5:pRR)zh p1me_ 7zQh1t7h ;RR):qRhaqz)pR2
RsRRCs0kMhRz)m 1p7e _1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMvQQhv5zvpa,Rmh_z1hQt )75,'RpDoCM02E2;R
RCRM8VOkM0MHFRhvQQvvz;R

RR--QR8:B.3c
VRRk0MOHRFMvQQhvRzv5:pRR)zh p1me_ 71hQt R7;)RR:Q hat2 )
RRRR0sCkRsMz h)1emp 17_Q th7#RH
LRRCMoH
RRRR0sCkRsMvQQhv5zvpa,RmQ_1t7h 5R),pC'DMEo02
2;RMRC8kRVMHO0FvMRQvhQz
v;
-RR-=R==========================================================================
=
R-R-R:Q8RcB3dR
RVOkM0MHFRXvqQvvzR,5pR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h R
H#RRRRO#FM00NMRZ1Q RR:hzqa)Rqp:v=RqvXQzpv5'MDCo,0ERD)'C0MoE
2;RRRRPHNsNCLDR4pjRRR:z h)1emp z7_ht1Qh5 71 QZ-84RF0IMF2Rj;R
RRNRPsLHND)CRjR4R:hRz)m 1p7e _1zhQ th7Q51Z4 -RI8FMR0Fj
2;RCRLo
HMRRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CsMRCs0kMqRhzR;
RCRRMH8RVR;
RpRRj:4R=mRa_5j4)Q 1Zp 5,QR1Z, 2R''X2R;
RHRRVpR5jp45jD4'C2V0R'=RXR'20MECR0sCkRsMp;j4
RRRR8CMR;HV
RRRR4)jRR:=ajm_4 5)1 QZ5R),1 QZ2',RX;'2
RRRRRHV54)j54)j'VDC0=2RR''X2ER0CsMRCs0kMjR)4R;
RCRRMH8RVR;
RHRRVhRz1hQt p7_ 511p,j4R4)j2ER0CRM
RRRRR0sCkRsM);j4
RRRR#CDCR
RRRRRskC0spMRj
4;RRRRCRM8H
V;RMRC8kRVMHO0FvMRqvXQz
v;
-RR-8RQ:3RBcRc
RMVkOF0HMqRvXzQvvpR5,RR):hRz)m 1p7e _t1Qh2 7R0sCkRsMz h)1emp 17_Q th7#RH
RRRRMOF#M0N0QR1Z: RRahqzp)qRR:=vQqXv5zvpC'DMEo0,'R)DoCM0;E2
RRRRsPNHDNLCjRp4:RRR)zh p1me_ 71hQt 175Q-Z 4FR8IFM0R;j2
RRRRsPNHDNLCjR)4:RRR)zh p1me_ 71hQt 175Q-Z 4FR8IFM0R;j2
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RERCMskC0shMRq
1;RRRRCRM8H
V;RRRRpRj4:a=Rm4_j51) Q5Z p1,RQ2Z ,XR''
2;RRRRH5VRp5j4p'j4D0CV2RR='2X'RC0EMCRs0MksR4pj;R
RRMRC8VRH;R
RRjR)4=R:R_amj)45 Z1Q ,5)RZ1Q R2,'2X';R
RRVRHRj5)4j5)4C'DVR02=XR''02RERCMskC0s)MRj
4;RRRRCRM8H
V;RRRRH1VRQ th7 _p1p15jR4,)2j4RC0EMR
RRRRRskC0s)MRj
4;RRRRCCD#
RRRRsRRCs0kMjRp4R;
RCRRMH8RVR;
R8CMRMVkOF0HMqRvXzQvv
;
R-R-R:Q8RcB36R
RVOkM0MHFRXvqQvvzRR5p:qRhaqz)p);RRz:Rh1) m pe7h_z1hQt 
72RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksRXvqQvvz5_amzQh1t7h 5Rp,)C'DMEo02),R2R;
R8CMRMVkOF0HMqRvXzQvv
;
R-R-R:Q8RcB3nR
RVOkM0MHFRXvqQvvzRR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksRXvqQvvz5_am1hQt p75,'R)DoCM0,E2R;)2
CRRMV8Rk0MOHRFMvQqXv;zv
R
R-Q-R8B:R3
c(RkRVMHO0FvMRqvXQz5vRpRR:z h)1emp z7_ht1Qh; 7R:)RRahqzp)q2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0svMRqvXQzpv5,mRa_1zhQ th7,5)RDp'C0MoE;22
CRRMV8Rk0MOHRFMvQqXv;zv
R
R-Q-R8B:R3
cURkRVMHO0FvMRqvXQz5vRpRR:z h)1emp 17_Q th7);RRQ:Rhta  
)2RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0svMRqvXQzpv5,mRa_t1Qh5 7)p,R'MDCo20E2R;
R8CMRMVkOF0HMqRvXzQvv
;
R-R-R============================================================================R

RR--QR8:Bg3c
VRRk0MOHRFM""?>R,5pR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RHRRV5R5pC'DMEo0R4<R2sRFR'5)DoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRz"hvQ )Ba_17"3"?">":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRsVFRHHRM'RpsoNMCFRDFRb
RRRRRHRRV5RpH=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7">"?"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7">"?"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRRHVQX#_5Rp2FQsR#5_X)02RE
CMRRRRRRRRskC0s'MRX
';RRRRRDRC#RHVpRR>)ER0CRM
RRRRRsRRCs0kM4R''R;
RRRRR#CDCR
RRRRRRCRs0MksR''j;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;>"
R
R-Q-R8B:R3
6jRkRVMHO0F"MR?R>"5Rp,)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0hR"z)v Q1B_a"73""?>"M:RkRDD8CC0O80C,CRs0MksHRMoXR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRFRVsRRHHpMR'MsNoDCRF
FbRRRRRRRRHpVR5RH2=-R''ER0CRM
RRRRRRRRRbsCFRs0"vhz B)Q_71a3?"">:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s'MRX
';RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRFRVsRRHH)MR'MsNoDCRF
FbRRRRRRRRH)VR5RH2=-R''ER0CRM
RRRRRRRRRbsCFRs0"vhz B)Q_71a3?"">:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s'MRX
';RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRVRHR_Q#X25pRRFsQX#_5R)20MEC
RRRRRRRR0sCkRsM';X'
RRRRCRRDV#HR>pRR0)RE
CMRRRRRRRRskC0s'MR4
';RRRRRDRC#RC
RRRRRsRRCs0kMjR''R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:B436
VRRk0MOHRFM""?>RR5p:qRhaqz)p);RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMazm_ht1Qh5 7p),R'MDCo20ERR?>)R;
R8CMRMVkOF0HM?R">
";
-RR-8RQ:3RB6R.
RMVkOF0HM?R">5"RpRR:Q hat; )R:)RR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMa1m_Q th7,5pRD)'C0MoE?2R>;R)
CRRMV8Rk0MOHRFM""?>;R

RR--QR8:Bd36
VRRk0MOHRFM""?>RR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp>R?R_amzQh1t7h 5R),pC'DMEo02R;
R8CMRMVkOF0HM?R">
";
-RR-8RQ:3RB6Rc
RMVkOF0HM?R">5"RpRR:z h)1emp 17_Q th7);RRQ:Rhta  R)2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp>R?R_am1hQt )75,'RpDoCM0;E2
CRRMV8Rk0MOHRFM""?>;R

RR--============================================================================
R
R-Q-R8B:R3
66RkRVMHO0F"MR?R<"5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0"vhz B)Q_71a3?""<:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRVRFsHMRHRsp'NCMoRFDFbR
RRRRRRVRHRHp52RR='R-'0MEC
RRRRRRRRsRRCsbF0hR"z)v Q1B_a"73""?<"':R-V'RF8kMRRHMObFlNRsC#H0sM
o"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0MksR''X;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRVRFsHMRHRs)'NCMoRFDFbR
RRRRRRVRHRH)52RR='R-'0MEC
RRRRRRRRsRRCsbF0hR"z)v Q1B_a"73""?<"':R-V'RF8kMRRHMObFlNRsC#H0sM
o"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0MksR''X;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRHQVR#5_XpF2Rs#RQ_)X52ER0CRM
RRRRRsRRCs0kMXR''R;
RRRRR#CDHpVRR)<RRC0EMR
RRRRRRCRs0MksR''4;R
RRRRRCCD#
RRRRRRRR0sCkRsM';j'
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
-RR-8RQ:3RB6Rn
RMVkOF0HM?R"<5"Rp),RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RHRRV5R5pC'DMEo0R4<R2sRFR'5)DoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRz"hvQ )Ba_17"3"?"<":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRsVFRHHRM'RpsoNMCFRDFRb
RRRRRHRRV5RpH=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7"<"?"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7"<"?"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRRHVQX#_5Rp2FQsR#5_X)02RE
CMRRRRRRRRskC0s'MRX
';RRRRRDRC#RHVpRR<)ER0CRM
RRRRRsRRCs0kM4R''R;
RRRRR#CDCR
RRRRRRCRs0MksR''j;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
6(RkRVMHO0F"MR?R<"5:pRRahqzp)q;RR):hRz)m 1p7e _1zhQ th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0saMRmh_z1hQt p75,'R)DoCM0RE2?)<R;R
RCRM8VOkM0MHFR<"?"
;
R-R-R:Q8R6B3UR
RVOkM0MHFR<"?"pR5RQ:Rhta  R);)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0saMRmQ_1t7h 5Rp,)C'DMEo02<R?R
);RMRC8kRVMHO0F"MR?;<"
R
R-Q-R8B:R3
6gRkRVMHO0F"MR?R<"5:pRR)zh p1me_ 7zQh1t7h ;RR):qRhaqz)ps2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0spMRRR?<azm_ht1Qh5 7)p,R'MDCo20E;R
RCRM8VOkM0MHFR<"?"
;
R-R-R:Q8RnB3jR
RVOkM0MHFR<"?"pR5Rz:Rh1) m pe7Q_1t7h ;RR):hRQa  t)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0spMRRR?<a1m_Q th7,5)RDp'C0MoE
2;RMRC8kRVMHO0F"MR?;<"
R
R-=-R=========================================================================
==
-RR-8RQ:3RBnR4
RMVkOF0HM?R"<R="5Rp,)RR:z h)1emp z7_ht1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0"vhz B)Q_71a3?""<"=":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRsVFRHHRM'RpsoNMCFRDFRb
RRRRRHRRV5RpH=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7"<"?=:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s'MRX
';RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRFRVsRRHH)MR'MsNoDCRF
FbRRRRRRRRH)VR5RH2=-R''ER0CRM
RRRRRRRRRbsCFRs0"vhz B)Q_71a3?""<"=":-R''FRVkRM8HOMRFNlbs#CR0MsHoR"
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCkRsM';X'
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRHRRV#RQ_pX52sRFR_Q#X25)RC0EMR
RRRRRRCRs0MksR''X;R
RRRRRCHD#VRRp<)=RRC0EMR
RRRRRRCRs0MksR''4;R
RRRRRCCD#
RRRRRRRR0sCkRsM';j'
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
n.RkRVMHO0F"MR?"<=R,5pR:)RR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbs"0Rh zv)_QB13a7"<"?=:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRVRFsHMRHRsp'NCMoRFDFbR
RRRRRRVRHRHp52RR='R-'0MEC
RRRRRRRRsRRCsbF0hR"z)v Q1B_a"73"=?<"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7"<"?=:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s'MRX
';RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRVRHR_Q#X25pRRFsQX#_5R)20MEC
RRRRRRRR0sCkRsM';X'
RRRRCRRDV#HR<pR=RR)0MEC
RRRRRRRR0sCkRsM';4'
RRRRCRRD
#CRRRRRRRRskC0s'MRj
';RRRRRMRC8VRH;R
RRMRC8VRH;R
RCRM8VOkM0MHFR<"?=
";
-RR-8RQ:3RBnRd
RMVkOF0HM?R"<R="5:pRRahqzp)q;RR):hRz)m 1p7e _1zhQ th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0saMRmh_z1hQt p75,'R)DoCM0RE2?R<=)R;
R8CMRMVkOF0HM?R"<;="
R
R-Q-R8B:R3
ncRkRVMHO0F"MR?"<=RR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMmRa_t1Qh5 7p),R'MDCo20ER=?<R
);RMRC8kRVMHO0F"MR?"<=;R

RR--QR8:B63n
VRRk0MOHRFM"=?<"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:hzqa)2qpR0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR?pR<a=Rmh_z1hQt )75,'RpDoCM0;E2
CRRMV8Rk0MOHRFM"=?<"
;
R-R-R:Q8RnB3nR
RVOkM0MHFR<"?=5"RpRR:z h)1emp 17_Q th7);RRQ:Rhta  R)2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp<R?=mRa_t1Qh5 7)p,R'MDCo20E;R
RCRM8VOkM0MHFR<"?=
";
-RR-=R==========================================================================
=
R-R-R:Q8RnB3(R
RVOkM0MHFR>"?=5"Rp),RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbs"0Rh zv)_QB13a7">"?=:""RDMkDCR800COCR8,skC0sMMHo"RX
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsM';X'
RRRR#CDCR
RRRRRVRFsHMRHRsp'NCMoRFDFbR
RRRRRRVRHRHp52RR='R-'0MEC
RRRRRRRRsRRCsbF0hR"z)v Q1B_a"73"=?>"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRsFCbs"0Rh zv)_QB13a7">"?=:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s'MRX
';RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRVRHR_Q#X25pRRFsQX#_5R)20MEC
RRRRRRRR0sCkRsM';X'
RRRRCRRDV#HR>pR=RR)0MEC
RRRRRRRR0sCkRsM';4'
RRRRCRRD
#CRRRRRRRRskC0s'MRj
';RRRRRMRC8VRH;R
RRMRC8VRH;R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RBnRU
RMVkOF0HM?R">R="5Rp,)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0hR"z)v Q1B_a"73"=?>"R":MDkDR08CCCO08s,RCs0kMoHMR
X"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s'MRX
';RRRRCCD#
RRRRVRRFHsRRRHMpN'sMRoCDbFF
RRRRRRRRRHVp25HR'=R-0'RE
CMRRRRRRRRRCRsb0FsRz"hvQ )Ba_17"3"?">="':R-V'RF8kMRRHMObFlNRsC#H0sM
o"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0MksR''X;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRVRFsHMRHRs)'NCMoRFDFbR
RRRRRRVRHRH)52RR='R-'0MEC
RRRRRRRRsRRCsbF0hR"z)v Q1B_a"73"=?>"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMXR''R;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRRHVQX#_5Rp2FQsR#5_X)02RE
CMRRRRRRRRskC0s'MRX
';RRRRRDRC#RHVp=R>R0)RE
CMRRRRRRRRskC0s'MR4
';RRRRRDRC#RC
RRRRRsRRCs0kMjR''R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?>"
;
R-R-R:Q8RnB3gR
RVOkM0MHFR>"?=5"RpRR:hzqa);qpR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMmRa_1zhQ th7,5pRD)'C0MoE?2R>)=R;R
RCRM8VOkM0MHFR>"?=
";
-RR-8RQ:3RB(Rj
RMVkOF0HM?R">R="5:pRRaQh )t ;RR):hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR_am1hQt p75,'R)DoCM0RE2?R>=)R;
R8CMRMVkOF0HM?R">;="
R
R-Q-R8B:R3
(4RkRVMHO0F"MR?">=RR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp>R?=mRa_1zhQ th7,5)RDp'C0MoE
2;RMRC8kRVMHO0F"MR?">=;R

RR--QR8:B.3(
VRRk0MOHRFM"=?>"pR5Rz:Rh1) m pe7Q_1t7h ;RR):hRQa  t)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0spMRR=?>R_am1hQt )75,'RpDoCM0;E2
CRRMV8Rk0MOHRFM"=?>"
;
R-R-R============================================================================R

RR--QR8:Bd3(
VRRk0MOHRFM""?=R,5pR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0p _pwRaRRRRRRRRR:hRQa  t)=R:RDp'C0MoE;-4
RRRRMOF#M0N0_R)pa wRRRRRRRRRRR:Q hatR ):)=R'MDCo-0E4R;
RNRRD#HNRRXpRRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7_5ppa wRI8FMR0FjH2R#;Rp
RRRRHNDNX#R)RRRRRRRRRRRRRRRRRR:z h)1emp z7_ht1Qh5 7) _pw8aRF0IMF2RjRRH#)R;
RORRF0M#NRM01 QZRRRRRRRRRRRR:qRhaqz)p=R:RXvqQvvz5Dp'C0MoE),R'MDCo20E;R
RRNRPsLHNDpCRXRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h 5Z1Q R-48MFI0jFR2R;
RPRRNNsHLRDC)RXRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7Q51Z4 -RI8FMR0Fj
2;RRRRPHNsNCLDR#sCk,D0R#sCk4D0R1:Raz7_pQmtBR;R-s-RCD#k0R
RLHCoMR
RR-R-RopFHDONDH$R80CMHDONRR0FN"MR=F"RbNCs03Fs
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbs"0Rh zv)_QB13a7"="?"R":MDkDR08CCCO08s,RCs0kMoHMR
X"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s'MRX
';RRRRCCD#
RRRRpRRXRRRR=R:R1) Q5Z XRp,1 QZ2R;
RRRRRR)XRRRR:)=R Z1Q )5X,QR1Z; 2
RRRRsRRCD#k0=R:R''4;R
RRRRRVRFsHMRHR'pXDRFI0pFRXH'EoDERF
FbRRRRRRRRskC#DR04:p=RX25HRR?=)HX52R;
RRRRRHRRVCRs#0kD4RR='Rz'0MEC
RRRRRRRRsRRCs0kMzR''R;
RRRRRCRRDV#HR#sCk4D0R'=RXF'RsCRs#0kDR'=RX0'RE
CMRRRRRRRRRCRs#0kDRR:=';X'
RRRRRRRR#CDCR
RRRRRRRRRskC#D:0R=CRs#0kDR8NMR#sCk4D0;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(Rc
RMVkOF0HM?R"=5"Rp),RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0p _pwRaRRRRRRRRR:hRQa  t)=R:RDp'C0MoE;-4
RRRRMOF#M0N0_R)pa wRRRRRRRRRRR:Q hatR ):)=R'MDCo-0E4R;
RNRRD#HNRRXpRRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh5 7p _pw8aRF0IMF2RjRRH#pR;
RNRRD#HNRRX)RRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh5 7) _pw8aRF0IMF2RjRRH#)R;
RORRF0M#NRM01 QZRRRRRRRRRRRR:qRhaqz)p=R:RXvqQvvz5Dp'C0MoE),R'MDCo20E;R
RRNRPsLHNDpCRXRRRRRRRRRRRR:RRR)zh p1me_ 71hQt 175Q-Z 4FR8IFM0R;j2
RRRRsPNHDNLCXR)RRRRRRRRRRRRRRR:z h)1emp 17_Q th7Q51Z4 -RI8FMR0Fj
2;RRRRPHNsNCLDR#sCk,D0R#sCk4D0R1:Raz7_pQmtBR;R-s-RCD#k0R
RLHCoM-RR-=R?
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbs"0Rh zv)_QB13a7"="?"R":MDkDR08CCCO08s,RCs0kMoHMR
X"RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRskC0s'MRX
';RRRRCCD#
RRRRpRRXRRRR=R:R1) Q5Z XRp,1 QZ2R;
RRRRRR)XRRRR:)=R Z1Q )5X,QR1Z; 2
RRRRsRRCD#k0=R:R''4;R
RRRRRVRFsHMRHR'pXDRFI0pFRXH'EoDERF
FbRRRRRRRRskC#DR04:p=RX25HRR?=)HX52R;
RRRRRHRRVCRs#0kD4RR='Rz'0MEC
RRRRRRRRsRRCs0kMzR''R;
RRRRRCRRDV#HR#sCk4D0R'=RXF'RsCRs#0kDR'=RX0'RE
CMRRRRRRRRRCRs#0kDRR:=';X'
RRRRRRRR#CDCR
RRRRRRRRRskC#D:0R=CRs#0kDR8NMR#sCk4D0;R
RRRRRRMRC8VRH;R
RRRRRCRM8DbFF;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(R6
RMVkOF0HM?R"=5"RpRR:hzqa);qpR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMmRa_1zhQ th7,5pRD)'C0MoE?2R=;R)
CRRMV8Rk0MOHRFM""?=;R

RR--QR8:Bn3(
VRRk0MOHRFM""?=RR5p:hRQa  t));RRz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMmRa_t1Qh5 7p),R'MDCo20ERR?=)R;
R8CMRMVkOF0HM?R"=
";
-RR-8RQ:3RB(R(
RMVkOF0HM?R"=5"RpRR:z h)1emp z7_ht1Qh; 7R:)RRahqzp)q2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMRRp?a=Rmh_z1hQt )75,'RpDoCM0;E2
CRRMV8Rk0MOHRFM""?=;R

RR--QR8:BU3(
VRRk0MOHRFM""?=RR5p:hRz)m 1p7e _t1Qh; 7R:)RRaQh )t 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMRRp?a=RmQ_1t7h 5R),pC'DMEo02R;
R8CMRMVkOF0HM?R"=
";
-RR-=R==========================================================================
=
R-R-R:Q8R(B3gR
RVOkM0MHFR/"?=5"Rp),RRz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0_Rppa wRRRRRRRRRRR:Q hatR ):p=R'MDCo-0E4R;
RORRF0M#NRM0) _pwRaRRRRRRRRR:hRQa  t)=R:RD)'C0MoE;-4
RRRRHNDNX#RpRRRRRRRRRRRRRRRRRR:z h)1emp z7_ht1Qh5 7p _pw8aRF0IMF2RjRRH#pR;
RNRRD#HNRRX)RRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7_5)pa wRI8FMR0FjH2R#;R)
RRRRMOF#M0N0QR1ZR RRRRRRRRRRRR:hzqa)Rqp:v=RqvXQzpv5'MDCo,0ERD)'C0MoE
2;RRRRPHNsNCLDRRpXRRRRRRRRRRRRRz:Rh1) m pe7h_z1hQt 175Q-Z 4FR8IFM0R;j2
RRRRsPNHDNLCXR)RRRRRRRRRRRRRRR:z h)1emp z7_ht1Qh5 71 QZ-84RF0IMF2Rj;R
RRNRPsLHNDsCRCD#k0s,RCD#k0:4RR71a_mzpt;QBR-R-R#sCk
D0RCRLoRHMRR--?R=
RHRRV5R5pC'DMEo0R4<R2sRFR'5)DoCM0<ERR242RC0EMR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRz"hvQ )Ba_17"3"?"/="M:RkRDD8CC0O80C,CRs0MksHRMoXR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRXRpRRRRRR:=)Q 1ZX 5p1,RQ2Z ;R
RRRRR)RXRR:RR= R)1 QZ5,X)RZ1Q 
2;RRRRRCRs#0kDRR:=';j'
RRRRVRRFHsRRRHMpDX'F0IRFXRp'oEHEFRDFRb
RRRRRsRRCD#k0:4R=XRp5RH2?R/=)HX52R;
RRRRRHRRVCRs#0kD4RR='Rz'0MEC
RRRRRRRRsRRCs0kMzR''R;
RRRRRCRRDV#HR#sCk4D0R'=RXF'RsCRs#0kDR'=RX0'RE
CMRRRRRRRRRCRs#0kDRR:=';X'
RRRRRRRR#CDCR
RRRRRRRRRskC#D:0R=CRs#0kDRRFsskC#D;04
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR/"?=
";
-RR-8RQ:3RBURj
RMVkOF0HM?R"/R="5Rp,)RR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRpp_ RwaRRRRRRRRRQ:Rhta  :)R='RpDoCM04E-;R
RRFROMN#0M)0R_wp aRRRRRRRR:RRRaQh )t RR:=)C'DMEo0-
4;RRRRNNDH#pRXRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h 5pp_ Rwa8MFI0jFR2#RHR
p;RRRRNNDH#)RXRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h 5p)_ Rwa8MFI0jFR2#RHR
);RRRRO#FM00NMRZ1Q RRRRRRRRRRRRh:Rq)azq:pR=qRvXzQvv'5pDoCM0RE,)C'DMEo02R;
RPRRNNsHLRDCpRXRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh5 71 QZ-84RF0IMF2Rj;R
RRNRPsLHND)CRXRRRRRRRRRRRR:RRR)zh p1me_ 71hQt 175Q-Z 4FR8IFM0R;j2
RRRRsPNHDNLCCRs#0kD,CRs#0kD4RR:1_a7ztpmQRB;RR--skC#DR0
RoLCHRMR-?-R=R
RRVRHRp55'MDCoR0E<2R4RRFs5D)'C0MoERR<4R220MEC
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0"vhz B)Q_71a3?""/"=":kRMD8DRCO0C0,C8R0sCkHsMMXoR"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRRpXRRRR:)=R Z1Q p5X,QR1Z; 2
RRRR)RRXRRRR=R:R1) Q5Z XR),1 QZ2R;
RRRRR#sCkRD0:'=Rj
';RRRRRFRVsRRHHpMRXF'DIFR0R'pXEEHoRFDFbR
RRRRRRCRs#0kD4=R:R5pXH?2R/)=RX25H;R
RRRRRRVRHR#sCk4D0R'=Rz0'RE
CMRRRRRRRRRCRs0MksR''z;R
RRRRRRDRC#RHVskC#DR04=XR''sRFR#sCkRD0=XR''ER0CRM
RRRRRRRRR#sCkRD0:'=RX
';RRRRRRRRCCD#
RRRRRRRRsRRCD#k0=R:R#sCkRD0FssRCD#k0
4;RRRRRRRRCRM8H
V;RRRRRMRC8FRDF
b;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?/"
;
R-R-R:Q8RUB34R
RVOkM0MHFR/"?=5"RpRR:hzqa);qpR:)RR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMmRa_1zhQ th7,5pRD)'C0MoE?2R/)=R;R
RCRM8VOkM0MHFR/"?=
";
-RR-8RQ:3RBUR.
RMVkOF0HM?R"/R="5:pRRaQh )t ;RR):hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksR_am1hQt p75,'R)DoCM0RE2?R/=)R;
R8CMRMVkOF0HM?R"/;="
R
R-Q-R8B:R3
UdRkRVMHO0F"MR?"/=RR5p:hRz)m 1p7e _1zhQ th7);RRh:Rq)azqRp2skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMp/R?=mRa_1zhQ th7,5)RDp'C0MoE
2;RMRC8kRVMHO0F"MR?"/=;R

RR--QR8:Bc3U
VRRk0MOHRFM"=?/"pR5Rz:Rh1) m pe7Q_1t7h ;RR):hRQa  t)s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0spMRR=?/R_am1hQt )75,'RpDoCM0;E2
CRRMV8Rk0MOHRFM"=?/"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413(#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14R(
RMVkOF0HM#R"DRN"5tq)Rz:Rh1) m pe7h_z1hQt R7;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp z7_ht1QhR 7HR#
RoLCHRM
RHRRVBR5mazhRR>=j02RE
CMRRRRRCRs0MksRQ1]wpa_ 5waq,)tRzBmh;a2
RRRR#CDCR
RRRRRskC0s1MR]aQw_t)Q]qa5)Rt,-zBmh;a2
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"N#D"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413U#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14RU
RMVkOF0HM#R"DRN"5tq)Rz:Rh1) m pe7Q_1t7h ;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _t1QhR 7HR#
RoLCHRM
RHRRVBR5mazhRR>=j02RE
CMRRRRRCRs0MksRQ1]wpa_ 5waq,)tRzBmh;a2
RRRR#CDCR
RRRRRskC0s1MR]aQw_t)Q]qa5)Rt,-zBmh;a2
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"N#D"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR413g#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R14Rg
RMVkOF0HM#R"sRN"5tq)Rz:Rh1) m pe7h_z1hQt R7;BhmzaRR:Q hat2 )
RRRR0sCkRsMz h)1emp z7_ht1QhR 7HR#
RoLCHRM
RHRRVBR5mazhRR>=j02RE
CMRRRRRCRs0MksRQ1]w)a_Qat]5tq),mRBz2ha;R
RRDRC#RC
RRRRR0sCkRsM1w]Qa _pwqa5)Rt,-zBmh;a2
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"N#s"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFR.13j#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3R1.Rj
RMVkOF0HM#R"sRN"5tq)Rz:Rh1) m pe7Q_1t7h ;mRBzRha:hRQa  t)R2
RsRRCs0kMhRz)m 1p7e _t1QhR 7HR#
RoLCHRM
RHRRVBR5mazhRR>=j02RE
CMRRRRRCRs0MksRQ1]w)a_Qat]5tq),mRBz2ha;R
RRDRC#RC
RRRRR0sCkRsM1w]Qa _pwqa5)Rt,-zBmh;a2
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"N#s"
;
RkRVMHO0FaMRmh_z1hQt 57RqR)t:qRhaqz)p1;RQ_Z )R 1:hRz)m 1p7e _1zhQ th7R2
RsRRCs0kMhRz)m 1p7e _1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMazm_ht1QhR 75tq)R>R=Rtq),R
RRRRRRRRRRRRRRRRRRRRRRQR1Z= R>QR1Z) _ D1'C0MoE
2;RMRC8kRVMHO0FaMRmh_z1hQt 
7;
VRRk0MOHRFMa1m_Q th7qR5):tRRaQh )t ;QR1Z) _ :1RR)zh p1me_ 71hQt 
72RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0saMRmQ_1t7h R)5qt=RR>)RqtR,
RRRRRRRRRRRRRRRRRRRRRZ1Q >R=RZ1Q  _)1C'DMEo02R;
R8CMRMVkOF0HMmRa_t1Qh; 7

RRRkRVMHO0F)MR Z1Q qR5)Rt,1 QZ_1) Rz:Rh1) m pe7h_z1hQt 
72RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR1) QRZ 5tq)RRRRR>R=Rtq),R
RRRRRRRRRRRRRRRRRRWh _Z1Q >R=RZ1Q  _)1C'DMEo02R;
R8CMRMVkOF0HM R)1 QZ;R

RMVkOF0HM R)1 QZR)5qt1,RQ_Z )R 1:hRz)m 1p7e _t1Qh2 7
RRRR0sCkRsMz h)1emp 17_Q th7#RH
LRRCMoH
RRRR0sCkRsM)Q 1Z5 RqR)tRRRRRR=>q,)t
RRRRRRRRRRRRRRRRRRRh_ W1 QZRR=>1 QZ_1) 'MDCo20E;R
RCRM8VOkM0MHFR1) Q;Z 
R
R-Q-R8p:R3R46
VRRk0MOHRFM"8NM"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7h_z1hQt 
72RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h RR5pNRM81_a7ztpmQeB_ mBa)25)2R;
R8CMRMVkOF0HMNR"M;8"
R
R-Q-R8p:R3R4n
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h Ra517p_zmBtQ_Be a5m)pN2RM)8R2R;
R8CMRMVkOF0HMNR"M;8"
R
R-Q-R8p:R3R4(
VRRk0MOHRFM""FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _1zhQ th7R2
RsRRCs0kMhRz)m 1p7e _1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMz h)1emp z7_ht1QhR 75FpRsaR17p_zmBtQ_Be a5m));22
CRRMV8Rk0MOHRFM""Fs;R

RR--QR8:pU34RR
RVOkM0MHFRs"F"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h Ra517p_zmBtQ_Be a5m)pF2Rs2R);R
RCRM8VOkM0MHFRs"F"
;
R-R-R:Q8R4p3gRR
RMVkOF0HMMR"N"M8RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _1zhQ th7R2
RsRRCs0kMhRz)m 1p7e _1zhQ th7#RH
LRRCMoH
RRRR0sCkRsMz h)1emp z7_ht1QhR 75MpRNRM81_a7ztpmQeB_ mBa)25)2R;
R8CMRMVkOF0HMMR"N"M8;R

RR--QR8:pj3.RR
RVOkM0MHFRN"MMR8"5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7h_z1hQt 57R1_a7ztpmQeB_ mBa)25pRMMN82R);R
RCRM8VOkM0MHFRN"MM;8"
R
R-Q-R8p:R3R.4
VRRk0MOHRFM"sMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7h_z1hQt 
72RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h RR5pMRFs1_a7ztpmQeB_ mBa)25)2R;
R8CMRMVkOF0HMMR"F;s"
R
R-Q-R8p:R3R..
VRRk0MOHRFM"sMF"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h Ra517p_zmBtQ_Be a5m)pM2RF)sR2R;
R8CMRMVkOF0HMMR"F;s"
R
R-Q-R8p:R3R.d
VRRk0MOHRFM"sGF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7h_z1hQt 
72RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h RR5pGRFs1_a7ztpmQeB_ mBa)25)2R;
R8CMRMVkOF0HMGR"F;s"
R
R-Q-R8p:R3R.c
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7h_z1hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h Ra517p_zmBtQ_Be a5m)pG2RF)sR2R;
R8CMRMVkOF0HMGR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3R.6HM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:p63.RR
RVOkM0MHFRM"GFRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 7zQh1t7h 2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7h_z1hQt 57RpMRGF1sRaz7_pQmtB _eB)am52)2;R
RCRM8VOkM0MHFRM"GF;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3R.nHM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:pn3.RR
RVOkM0MHFRM"GFRs"5:pRR)zh p1me_ 7zQh1t7h ;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7h_z1hQt 57R1_a7ztpmQeB_ mBa)25pRFGMs2R);R
RCRM8VOkM0MHFRM"GF;s"
R
R-Q-R8p:R3R.(
VRRk0MOHRFM"8NM"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt 57RpMRN8aR17p_zmBtQ_Be a5m));22
CRRMV8Rk0MOHRFM"8NM"
;
R-R-R:Q8R.p3URR
RMVkOF0HMNR"MR8"5:pRR)zh p1me_ 71hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h Ra517p_zmBtQ_Be a5m)pN2RM)8R2R;
R8CMRMVkOF0HMNR"M;8"
R
R-Q-R8p:R3R.g
VRRk0MOHRFM""FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _t1Qh2 7
RRRR0sCkRsMz h)1emp 17_Q th7#RH
LRRCMoH
RRRR0sCkRsMz h)1emp 17_Q th7pR5RRFs1_a7ztpmQeB_ mBa)25)2R;
R8CMRMVkOF0HMFR"s
";
-RR-8RQ:3Rpd
jRRkRVMHO0F"MRFRs"5:pRR)zh p1me_ 71hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h Ra517p_zmBtQ_Be a5m)pF2Rs2R);R
RCRM8VOkM0MHFRs"F"
;
R-R-R:Q8Rdp34RR
RMVkOF0HMMR"N"M8RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _t1Qh2 7
RRRR0sCkRsMz h)1emp 17_Q th7#RH
LRRCMoH
RRRR0sCkRsMz h)1emp 17_Q th7pR5RMMN8aR17p_zmBtQ_Be a5m));22
CRRMV8Rk0MOHRFM"MMN8
";
-RR-8RQ:3Rpd
.RRkRVMHO0F"MRM8NM"pR5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt 57R1_a7ztpmQeB_ mBa)25pRMMN82R);R
RCRM8VOkM0MHFRN"MM;8"
R
R-Q-R8p:R3Rdd
VRRk0MOHRFM"sMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt 57RpFRMsaR17p_zmBtQ_Be a5m));22
CRRMV8Rk0MOHRFM"sMF"
;
R-R-R:Q8Rdp3cRR
RMVkOF0HMMR"FRs"5:pRR)zh p1me_ 71hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h Ra517p_zmBtQ_Be a5m)pM2RF)sR2R;
R8CMRMVkOF0HMMR"F;s"
R
R-Q-R8p:R3Rd6
VRRk0MOHRFM"sGF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7Q_1t7h 2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt 57RpFRGsaR17p_zmBtQ_Be a5m));22
CRRMV8Rk0MOHRFM"sGF"
;
R-R-R:Q8Rdp3nRR
RMVkOF0HMGR"FRs"5:pRR)zh p1me_ 71hQt R7;)RR:1_a7ztpmQ
B2RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h Ra517p_zmBtQ_Be a5m)pG2RF)sR2R;
R8CMRMVkOF0HMGR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3Rd(HM#RFO0RFNlb0DHLCHRI0QER R  1R084nj(-U4g(B3RFCllMR0
RR--FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2VRFsQ   R810R(4jng-4UO(RFNlb0HHLD$H03R
R-----------------------------------------------------------------------------R-
RR--QR8:p(3dRR
RVOkM0MHFRM"GFRs"5:pRR71a_mzpt;QBR:)RR)zh p1me_ 71hQt 
72RRRRskC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h RR5pGsMFR71a_mzpt_QBea Bm))52
2;RMRC8kRVMHO0F"MRGsMF"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRdp3U#RHR0MFRlOFbHN0LRDCIEH0R Q  0R18jR4(4n-g3U(RlBFl0CM
-RR-kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVs RQ 1 R048Rj-(n4(gURlOFbHN0LHHD0
$3R-R-----------------------------------------------------------------------------
-RR-8RQ:3Rpd
URRkRVMHO0F"MRGsMF"pR5Rz:Rh1) m pe7Q_1t7h ;RR):aR17p_zmBtQ2R
RRCRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt 57R1_a7ztpmQeB_ mBa)25pRFGMs2R);R
RCRM8VOkM0MHFRM"GF;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RdgHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pg3d
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMMRN81R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMNR"M;8"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RcjHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pj3c
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMNRM8571a_mzpt_QBea Bm5)Rp;22
CRRMV8Rk0MOHRFM"8NM"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp34#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcR4
RMVkOF0HMMR"N"M8RR5p:hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRMMN81R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMMR"N"M8;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMp.3cRRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8Rcp3.R
RVOkM0MHFRN"MMR8"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMNRMM58R1_a7ztpmQeB_ mBa)pR52
2;RMRC8kRVMHO0F"MRM8NM"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3d#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcRd
RMVkOF0HMFR"s5"RpRR:z h)1emp 17_Q th7s2RCs0kMaR17p_zmBtQR
H#RCRLo
HMRRRRskC0sFMRs1R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMFR"s
";
-RR-----------------------------------------------------------------------------R
R-h-RF:0CRMwkOF0HM3RpcHcR#FRM0FROl0bNHCLDR0IHE8RCHF0HMF#RV RQ 1 R048RjR(nVlsF
-RR-gR4U0(REksFo.ERj3j.RlBFl0CMR0FkRC0ERMVkOF0HM8R5CNODsHN0FNMRML8RF28$RsVF
-RR-FROl0bNHDLHHR0$IEH0RC0E#CCR8HH0F3M#
-RR-----------------------------------------------------------------------------R
R-Q-R8p:R3
ccRkRVMHO0F"MRFRs"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMsRFRa517p_zmBtQ_Be aRm)52p2;R
RCRM8VOkM0MHFRs"F"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp36#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcR6
RMVkOF0HMMR"FRs"5:pRR)zh p1me_ 71hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMMRFs571a_mzpt_QBea Bm5)Rp;22
CRRMV8Rk0MOHRFM"sMF"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3n#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcRn
RMVkOF0HMMR"FRs"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMFRMs1R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMMR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3Rc(HM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:p(3c
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7Q_1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMFRGs1R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMGR"F;s"
R
R-----------------------------------------------------------------------------R-
RR--hCF0:kRwMHO0FpMR3RcUHM#RFO0RFNlb0DHLCHRI0CER8HH0FRM#FQVR R  1R084nj(RFVslR
R-4-RgRU(0FEskRoE..jj3FRBlMlC0kRF0ER0CkRVMHO0F5MR8DCON0sNHRFMNRM8L$F82FRVsR
R-O-RFNlb0HHLD$H0R0IHEER0CR#CC08HH#FM3R
R-----------------------------------------------------------------------------R-
RR--QR8:pU3c
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7h_z1hQt R72skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMGRFs571a_mzpt_QBea Bm5)Rp;22
CRRMV8Rk0MOHRFM"sGF"
;
R-R-----------------------------------------------------------------------------
-RR-FRh0RC:wOkM0MHFRcp3g#RHR0MFRlOFbHN0LRDCIEH0RHC80MHF#VRFR Q  0R18jR4(VnRs
FlR-R-RU4g(ER0soFkEjR.jR.3BlFlCRM0FRk00RECVOkM0MHFRC58OsDNNF0HMMRN8FRL8R$2V
FsR-R-RlOFbHN0LHHD0I$RHR0E0#ECC8RCHF0HM
#3R-R-----------------------------------------------------------------------------
-RR-8RQ:3RpcRg
RMVkOF0HMGR"M"FsRR5p:hRz)m 1p7e _t1Qh2 7R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRFGMs1R5az7_pQmtB _eB)amR25p2R;
R8CMRMVkOF0HMGR"M"Fs;R

R----------------------------------------------------------------------------
--R-R-R0hFCw:Rk0MOHRFMpj36RRH#MRF0ObFlNL0HDICRHR0EC08HH#FMRRFVQ   R810R(4jnsRVFRl
RR--4(gURs0EFEkoRj.j.B3RFCllMF0Rk00REVCRk0MOHRFM5O8CDNNs0MHFR8NMR8LF$V2RFRs
RR--ObFlNL0HH0DH$HRI00ERECC#RHC80MHF#R3
R----------------------------------------------------------------------------
--R-R-R:Q8R6p3jR
RVOkM0MHFRM"GFRs"5:pRR)zh p1me_ 7zQh1t7h 2CRs0MksR71a_mzptRQBHR#
RoLCHRM
RsRRCs0kMMRGF5sR1_a7ztpmQeB_ mBa)pR52
2;RMRC8kRVMHO0F"MRGsMF"
;
R-R-R:Q8Rda3
VRRk0MOHRFMaXm_j54R1RR:z h)1emp z7_ht1Qh2 7R0sCkRsMz h)1emp z7_ht1QhR 7HR#
RoLCHRM
RsRRCs0kMhRz)m 1p7e _1zhQ th7m5a_4Xj571a_mzpt_QBea Bm1)52;22
CRRMV8Rk0MOHRFMaXm_j
4;
-RR-8RQ:3RacR
RVOkM0MHFR_amXRj45:1RR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h 5_amX5j41_a7ztpmQeB_ mBa)2512
2;RMRC8kRVMHO0FaMRmj_X4
;
R-R-R:Q8R6a3
VRRk0MOHRFMaXm_jR4Z5:1RR)zh p1me_ 7zQh1t7h 2CRs0MksR)zh p1me_ 7zQh1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7h_z1hQt a75mj_X41Z5az7_pQmtB _eB)am52122R;
R8CMRMVkOF0HMmRa_4XjZ
;
R-R-R:Q8Rna3
VRRk0MOHRFMaXm_jR4Z5:1RR)zh p1me_ 71hQt R72skC0szMRh1) m pe7Q_1t7h R
H#RCRLo
HMRRRRskC0szMRh1) m pe7Q_1t7h 5_amXZj4571a_mzpt_QBea Bm1)52;22
CRRMV8Rk0MOHRFMaXm_j;4Z
R
R-Q-R8a:R3R(
RMVkOF0HMmRa_jzX41R5Rz:Rh1) m pe7h_z1hQt R72skC0szMRh1) m pe7h_z1hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 7zQh1t7h 5_amz4Xj571a_mzpt_QBea Bm1)52;22
CRRMV8Rk0MOHRFMazm_X;j4
R
R-Q-R8a:R3RU
RMVkOF0HMmRa_jzX41R5Rz:Rh1) m pe7Q_1t7h 2CRs0MksR)zh p1me_ 71hQt H7R#R
RLHCoMR
RRCRs0MksR)zh p1me_ 71hQt a75mX_zj145az7_pQmtB _eB)am52122R;
R8CMRMVkOF0HMmRa_jzX4
;
R-R-R:Q8Rga3
VRRk0MOHRFMQX1_RR51:hRz)m 1p7e _1zhQ th7s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMQX1_571a_mzpt_QBea Bm1)52
2;RMRC8kRVMHO0FQMR1;_X
R
R-Q-R8a:R3
4jRkRVMHO0FQMR1R_X5:1RR)zh p1me_ 71hQt R72skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR_Q1Xa517p_zmBtQ_Be a5m)1;22
CRRMV8Rk0MOHRFMQX1_;R
R

RRRRRR-=-R=========================================================================
==R-R-Rs#0HRMoOPFMCHs#FNMRMI8RsCH0RCFbsHN0F
M#R-R-R============================================================================R
R
RRRRMVkOF0HMFR0_s#0HRMo5DPNkRCRR:RRRRHMz h)1emp z7_ht1Qh2 7R0sCkRsM1Qa)hHtR#R
RRDRNHRN#HDPNkRCRRRR:z h)1emp z7_ht1Qh5 74FR0RDPNkDC'C0MoEH2R#NRPD;kC
RRRRsPNHDNLCCRs#0kDR1:Rah)QtR540PFRNCDk'MDCo20E;L
SCMoH
RRRRRHVPkNDCC'DMEo0R4<RRC0EMR
RRRRRskC0shMRz
1;RRRRCCD#
RRRRVRRFHsRRRHMHDPNksC'NCMoRFDFbR
RRRRRRCRs#0kD5RH2:v=Re_pg0OF_E5NsHDeNkHC52
2;RRRRRMRC8FRDF
b;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_0MsHoR;
RR
RVOkM0MHFR_0F#H0sM5oRPkNDCRRRRRR:HzMRh1) m pe7Q_1t7h 2CRs0MksR)1aQRhtHR#
RNRRD#HNRNHPDRkCR:RRR)zh p1me_ 71hQt 475RR0FPkNDCC'DMEo02#RHRDPNk
C;RRRRPHNsNCLDR#sCkRD0:aR1)tQh504RFNRPD'kCDoCM0;E2
LRRCMoH
RRRRRHVPkNDCC'DMEo0R4<RRC0EMR
RRRRRskC0shMRz
1;RRRRCCD#
RRRRVRRFHsRRRHMHDPNksC'NCMoRFDFbR
RRRRRRCRs#0kD5RH2:v=Re_pg0OF_E5NsHDeNkHC52
2;RRRRRMRC8FRDF
b;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_0MsHoR;
RR
RVOkM0MHFR_0FFs#0HRMo5DPNk:CRR)zh p1me_ 7zQh1t7h 2CRs0MksR)1aQRhtHR#
RoLCHRM
RsRRCs0kMFR0_0F#soHM571a_mzpt_QBea Bm5)RPkNDC;22
CRRMV8Rk0MOHRFM0FF_#H0sM
o;
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:z h)1emp 17_Q th7s2RCs0kMaR1)tQhR
H#RRRRO#FM00NMR#sCk_D0DoCM0:ERRaQh )t RR:=5DPNkDC'C0MoE2+./
d;RRRRO#FM00NMR8bNRRRRRRRRR:RRR71a_mzpt_QBea Bm4)5RR0F5#sCk_D0DoCM0dE*RR-
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRPkNDCC'DMEo02R2
RRRRRR:=5EF0CRs#=P>RNCDkRN5PD'kCD0CV2R2;RR-- CG0M#8RHRoML
H0RCRLo
HMRRRRskC0s0MRF#_F0MsHoN5b8RR&1_a7ztpmQeB_ mBa)PR5NCDk2
2;RMRC8kRVMHO0F0MRF#_F0MsHo
;
RkRVMHO0F0MRF#_E0MsHoPR5NCDkRz:Rh1) m pe7h_z1hQt R72skC0s1MRah)Qt#RH
LRRCMoH
RRRR0sCkRsM0EF_#H0sM1o5az7_pQmtB _eB)amRN5PD2kC2R;
R8CMRMVkOF0HMFR0_0E#soHM;R

RMVkOF0HMFR0_0E#soHMRN5PDRkC:hRz)m 1p7e _t1Qh2 7R0sCkRsM1Qa)hHtR#R
RRFROMN#0Ms0RCD#k0C_DMEo0RQ:Rhta  :)R=PR5NCDk'MDCo+0Edc2/;R
RRFROMN#0Mb0RNR8RRRRRRRRRR1:Raz7_pQmtB _eB)am504RFsR5CD#k0C_DMEo0*-cR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNRPD'kCDoCM02E2
RRRR:RR=FR50sEC#>R=RDPNk5CRPkNDCC'DV202;-RR-GR 08CMRo#HMHRL0R
RLHCoMR
RRCRs0MksR_0FEs#0H5MobRN8&aR17p_zmBtQ_Be aRm)5DPNk2C2;R
RCRM8VOkM0MHFR_0FEs#0H;Mo
C

Mh8Rz)v Q1B_a
7;
