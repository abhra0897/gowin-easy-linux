--
@ER--B$FbsEHo0OR52gR4g-cRRj.jd$R1MHbDO$H0ROQM
R--fN]C8:CsR#//$DMbH0OH$N/lb/oIlbNbC/s#GHHDMDG/HoL/CsMCHoO/CoM_CsMCHsO/Nsl__PI3E48yR-f
--

----RpB p)RXq.vdXR47-----H
DLssN$CRHC
C;kR#CHCCC38#0_oDFH4O_43ncN;DD
Ck#RCHCC03#8F_Do_HO#MHoCN83D
D;DsHLNRs$k#MHH
l;kR#Ck#MHHPl3ObFlFMMC0N#3D
D;
0CMHR0$Xv)qd4.X7#RH
bRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRRRR7RRRR:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:jRRRHM#_08koDFH
O;RRRRRRRR7qu)4RR:H#MR0k8_DHFoOR;
RRRRR7RRu.)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqd:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:cRRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRqX)vXd.4
7;NEsOHO0C0CksRqX)vXd.4e7_RRFVXv)qd4.X7#RH
SRR#MHoNIDRCRj,I,C4Rj#F,FR#48,RFRj,8:F4R8#0_oDFH
O;LHCoM7
Su<mR=FR8jERIC5MR7qu)cRR='2j'R#CDCFR84S;
1Rum<#=RFIjRERCM5Rqc=jR''C2RDR#C#;F4
CSIj=R<RRW NRM850MFR2qc;I
SC<4R= RWR8NMR;qc
zRSjRR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRIjW,RBRpi=W>RB,piRm7uRR=>8,FjRm1uRR=>#2Fj;S
Rz:4RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR4,WiBpRR=>WiBp,uR7m>R=R48F,uR1m>R=R4#F2C;
MX8R)dqv.7X4_
e;
----B-R RppXv)qn4cX7-R--
--DsHLNRs$HCCC;#
kCCRHC#C30D8_FOoH_n44cD3NDk;
#HCRC3CC#_08DHFoOH_#o8MC3DND;H
DLssN$MRkHl#H;#
kCMRkHl#H3FPOlMbFC#M03DND;C

M00H$)RXqcvnXR47HR#
RsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRRqR6RRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:6RRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRqX)vXnc4
7;NEsOHO0C0CksRqX)vXnc4e7_RRFVXv)qn4cX7#RH
SRR#MHoNIDRCRj,I,C4R.IC,CRId#,RFRj,#,F4R.#F,FR#d8,RFRj,8,F4R.8F,FR8d#:R0D8_FOoH;C
Lo
HMSm7uRR<=Rj8FRCIEM7R5u6)qR'=RjN'RM78Ruc)qR'=RjR'2CCD#RS
S8RF4IMECRu57)Rq6=jR''MRN8uR7)Rqc=4R''C2RDR#C
8SSFI.RERCM5)7uq=6RR''4R8NMR)7uq=cRR''j2DRC#
CRSFS8dS;
1Rum<R=R#RFjIMECR65qR'=RjN'RMq8RcRR='2j'R#CDCSR
S4#FRCIEMqR56RR='Rj'NRM8q=cRR''42DRC#
CRSFS#.ERIC5MRq=6RR''4R8NMRRqc=jR''C2RDR#C
#SSF
d;SjICRR<=WN RM58RMRF0qR62NRM850MFR2qc;I
SC<4R= RWR8NMRF5M06Rq2MRN8cRq;I
SC<.R= RWR8NMRRq6NRM850MFR2qc;I
SC<dR= RWR8NMRRq6NRM8q
c;RjSzR):Rqnv4XR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>7q,Rj>R=R,qjRRq4=q>R4q,R.>R=R,q.RRqd=q>RdR,
S7SSuj)qRR=>7qu)j7,Ru4)qRR=>7qu)47,Ru.)qRR=>7qu).7,Rud)qRR=>7qu)d
,RSWSS >R=RjIC,BRWp=iR>BRWpRi,7Rum=8>RFRj,1Rum=#>RF;j2
zRS4RR:)4qvn7X4RR
RRRRRRRRRRRRRRFRbsl0RN5bR7>R=RR7,q=jR>jRq,4RqRR=>qR4,q=.R>.Rq,dRqRR=>q
d,RSSS7qu)j>R=R)7uqRj,7qu)4>R=R)7uqR4,7qu).>R=R)7uqR.,7qu)d>R=R)7uqRd,
SSSW= R>CRI4W,RBRpi=W>RB,piRm7uRR=>8,F4Rm1uRR=>#2F4;S
Rz:.RRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>,R7RRqj=q>Rjq,R4>R=R,q4RRq.=q>R.q,Rd>R=R,qd
SRSS)7uq=jR>uR7),qjR)7uq=4R>uR7),q4R)7uq=.R>uR7),q.R)7uq=dR>uR7),qdRS
SSRW =I>RCR.,WiBpRR=>WiBp,uR7m>R=R.8F,uR1m>R=R.#F2R;
SRzd:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=7>R,jRqRR=>qRj,q=4R>4Rq,.RqRR=>qR.,q=dR>dRq,S
RSuS7)Rqj=7>Ruj)q,uR7)Rq4=7>Ru4)q,uR7)Rq.=7>Ru.)q,uR7)Rqd=7>Rud)q,SR
S SWRR=>I,CdRpWBi>R=RpWBi7,Ru=mR>FR8d1,Ru=mR>FR#d
2;CRM8Xv)qn4cX7;_e
-
-

---1-RHDlbCqR)vHRI0#ERHDMoC7Rq71) 1FRVsFRL0sERCRN8NRM8I0sHC-
-RsaNoRC0:HRXDGHM

--
LDHs$NsRCHCCk;
#HCRC3CC#_08DHFoO4_4nNc3D
D;kR#CHCCC38#0_oDFH#O_HCoM8D3NDD;
HNLssk$RMHH#lk;
#kCRMHH#lO3PFFlbM0CM#D3NDC;
M00H$qR)v__)W#RH
CSoMHCsO
R5SRRRRlVNHRD$:0R#soHMRR:="MMFC
";SHSI8R0E:MRH0CCos=R:RR4;
NSS8I8sHE80RH:RMo0CC:sR=;RnRRRRRRRR-L-RHCoRMoFkEFRVsCR8b
0ESCS8bR0E:MRH0CCos=R:R;cU
8SSF_k0sRCo:FRLFNDCM=R:RDVN#RC;RRRRRR--ERN#Fbk0ks0RCSo
SM8H_osCRL:RFCFDN:MR=NRVD;#CRRRRRRRR-E-RN8#RNR0NHkMb0CRsoS
Ss8N8sC_soRR:LDFFCRNM:V=RNCD#;RRRR-RR-NRE#CRsNN8R8C8s#s#RCSo
S8IN8ss_C:oRRFLFDMCNR=R:RDVN#RCRRRRR-E-RNI#RsCH0R8N8s#C#RosC
2SS;b
SFRs05S
S7amz:kRF00R#8F_Do_HOP0COFIs5HE80-84RF0IMF2Rj;S
S)7q7)RR:H#MR0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2S;
Sh7QRRR:H#MR0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2S;
S7Wq7:)RRRHM#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0Fj
2;S SWRRR:H#MR0D8_FOoH;RRRRRRR-I-RsCH0RNCMLRDCVRFss
NlSpSBiRR:H#MR0D8_FOoH;RRRRRRR-O-RD	FORsVFRlsN,8RN8Rs,8
HMSBSmp:iRRRHM#_08DHFoORRRRRRR-F-RbO0RD	FORsVFR8I_F
k0S;S2
8CMR0CMHR0$)_qv);_W
-
-
R--w#Hs0lRHblDCCNM00MHFR#lk0CRLRDONDRC8NEsOj-
-
ONsECH0Os0kCDRLF_O	sRNlF)VRq)v__HWR#F
OlMbFCRM0Xv)qd4.X7RRRb0FsRR5
RRRRR7RRuRmRRF:Rk#0R0k8_DHFoOR;RRRRRRRR
RRRRR1RRuRmRRF:Rk#0R0k8_DHFoO
;
RRRRRRRRqRjRRRR:H#MR0k8_DHFoOR;
RRRRRqRR4RRRRH:RM0R#8D_kFOoH;R
RRRRRR.RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqdR:RRRRHM#_08koDFH
O;RRRRRRRRqRcRRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRRpWBi:RRRRHM#_08koDFHRO;RRRRR
RRRRRRRRRRWR RRRR:H#MR0k8_DHFoOR
RRRRRRR2;RM
C8FROlMbFC;M0
lOFbCFMMX0R)nqvc7X4RbRRFRs05R
RRRRRRuR7mRRR:kRF00R#8D_kFOoH;RRRRRRRRR
RRRRRRuR1mRRR:kRF00R#8D_kFOoH;R

RRRRRqRRjRRRRH:RM0R#8D_kFOoH;R
RRRRRR4RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq.R:RRRRHM#_08koDFH
O;RRRRRRRRqRdRRRR:H#MR0k8_DHFoOR;
RRRRRqRRcRRRRH:RM0R#8D_kFOoH;R
RRRRRR6RqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRR7RRu6)qRH:RM0R#8D_kFOoH;R
RRRRRRBRWpRiR:MRHR8#0_FkDo;HORRRRRRRR
RRRRRRRRRW R:RRRRHM#_08koDFHRO
RRRRR;R2RCR
MO8RFFlbM0CM;k
VMHO0FVMRk_MOH0MH5:LRRFLFDMCN2CRs0MksRs#0HRMoHL#
CMoH
HRRVLR52ER0CRM
RsRRCs0kM"5"2R;
R#CDCR
RRCRs0Mks5F"BkRD8MRF0HDlbCMlC0DRAFRO	)3qvRRQ#0RECs8CNR8N8s#C#RosCHC#0sRC8kM#HoER0CNR#lOCRD	FORRN#0REC)?qv"
2;RMRC8VRH;M
C8kRVMHO_M;H0
MVkOF0HMCRo0M_C8C_8b50E#CHxRH:RMo0CC;sRRb8C0:ERR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRMlH_x#HCRR:HCM0oRCs:j=R;C
Lo
HMRHRlMH_#x:CR=CR8b;0E
HRRV#R5HRxC<CR8b20ERC0EMR
RRHRlMH_#x:CR=HR#x
C;RMRC8VRH;R
RskC0slMRH#M_H;xC
8CMR0oC_8CM_b8C0
E;Ns00H0LkCCRoMNCs0_FssFCbs:0RRs#0H;Mo
0N0skHL0oCRCsMCNs0F_bsCFRs0FLVRD	FO_lsNRN:RsHOE00COkRsCHV#Rk_MOH0MH58sN8ss_C;o2
R--LHCoMDRLFRO	sRNlHDlbCMlC0HN0F#MRHNoMD0#
$RbCH_M0NNss$#RHRsNsN5$RjFR0RR62FHVRMo0CC
s;O#FM00NMR8IH0NE_s$sNRH:RMN0_s$sNRR:=5R4,.c,R,,RgR,4UR2dn;F
OMN#0M80RCEb0_sNsN:$RR0HM_sNsN:$R=4R5ncdU,4RUgR.,cnjg,jR.cRU,4cj.,4R6.
2;O#FM00NMRP8Hd:.RR0HMCsoCRR:=58IH04E-2n/d;F
OMN#0M80RHnP4RH:RMo0CC:sR=IR5HE80-/424
U;O#FM00NMRP8HURR:HCM0oRCs:5=RI0H8E2-4/
g;O#FM00NMRP8HcRR:HCM0oRCs:5=RI0H8E2-4/
c;O#FM00NMRP8H.RR:HCM0oRCs:5=RI0H8E2-4/
.;O#FM00NMRP8H4RR:HCM0oRCs:5=RI0H8E2-4/
4;
MOF#M0N0FRLFRD4:FRLFNDCM=R:RH58P>4RR;j2
MOF#M0N0FRLFRD.:FRLFNDCM=R:RH58P>.RR;j2
MOF#M0N0FRLFRDc:FRLFNDCM=R:RH58P>cRR;j2
MOF#M0N0FRLFRDU:FRLFNDCM=R:RH58P>URR;j2
MOF#M0N0FRLFnD4RL:RFCFDN:MR=8R5HnP4Rj>R2O;
F0M#NRM0LDFFd:.RRFLFDMCNRR:=5P8Hd>.RR;j2
F
OMN#0M80RHnP4dRUc:MRH0CCos=R:RC58b-0E442/ncdU;F
OMN#0M80RH4PUg:.RR0HMCsoCRR:=5b8C04E-24/Ug
.;O#FM00NMRP8HcnjgRH:RMo0CC:sR=8R5CEb0-/42cnjg;F
OMN#0M80RHjP.c:URR0HMCsoCRR:=5b8C04E-2j/.c
U;O#FM00NMRP8H4cj.RH:RMo0CC:sR=8R5CEb0-/424cj.;F
OMN#0M80RH4P6.RR:HCM0oRCs:5=R80CbE2-4/.64;O

F0M#NRM0LDFF6R4.:FRLFNDCM=R:RH58P.64Rj>R2O;
F0M#NRM0LDFF4cj.RL:RFCFDN:MR=8R5HjP4.>cRR;j2
MOF#M0N0FRLFjD.c:URRFLFDMCNRR:=5P8H.UjcRj>R2O;
F0M#NRM0LDFFcnjgRL:RFCFDN:MR=8R5HjPcg>nRR;j2
MOF#M0N0FRLF4DUg:.RRFLFDMCNRR:=5P8HU.4gRj>R2O;
F0M#NRM0LDFF4UndcRR:LDFFCRNM:5=R84HPncdURj>R2
;
O#FM00NMRl#k_8IH0:ERR0HMCsoCRR:=Apmm 'qhb5F#LDFF4+2RRmAmph q'#bF5FLFDR.2+mRAmqp hF'b#F5LF2DcRA+Rm mpqbh'FL#5FUFD2RR+Apmm 'qhb5F#LDFF4;n2
MOF#M0N0kR#lC_8bR0E:MRH0CCos=R:R-6RRm5Amqp hF'b#F5LF4D6.+2RRmAmph q'#bF5FLFD.4jc+2RRmAmph q'#bF5FLFDc.jU+2RRmAmph q'#bF5FLFDgcjn+2RRmAmph q'#bF5FLFDgU4.;22
F
OMN#0MI0R_FOEH_OCI0H8ERR:HCM0oRCs:I=RHE80_sNsN#$5kIl_HE802O;
F0M#NRM0IE_OFCHO_b8C0:ERR0HMCsoCRR:=80CbEs_Ns5N$#_klI0H8E
2;O#FM00NMRO8_EOFHCH_I8R0E:MRH0CCos=R:R8IH0NE_s$sN5l#k_b8C0;E2
MOF#M0N0_R8OHEFO8C_CEb0RH:RMo0CC:sR=CR8b_0ENNss$k5#lC_8b20E;O

F0M#NRM0IH_I8_0EM_klODCD#RR:HCM0oRCs:5=RI0H8E2-4/OI_EOFHCH_I8R0E+;R4
MOF#M0N0_RI80CbEk_MlC_ODRD#:MRH0CCos=R:RC58b-0E4I2/_FOEH_OC80CbERR+4
;
O#FM00NMRI8_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/8OHEFOIC_HE80R4+R;F
OMN#0M80R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/428E_OFCHO_b8C0+ERR
4;
MOF#M0N0_RI#CHxRH:RMo0CC:sR=_RII0H8Ek_MlC_ODRD#*_RI80CbEk_MlC_OD;D#
MOF#M0N0_R8#CHxRH:RMo0CC:sR=_R8I0H8Ek_MlC_ODRD#*_R880CbEk_MlC_OD;D#
F
OMN#0ML0RF_FD8RR:LDFFCRNM:5=R8H_#x-CRR#I_HRxC<j=R2O;
F0M#NRM0LDFF_:IRRFLFDMCNRR:=M5F0LDFF_;82
F
OMN#0MO0REOFHCH_I8R0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCH_I820E;F
OMN#0MO0REOFHCC_8bR0E:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_2RR*8E_OFCHO_b8C0RE2+AR5m mpqbh'FL#5F_FDI*2RROI_EOFHCC_8b20E;F
OMN#0MI0RHE80_lMk_DOCD:#RR0HMCsoCRR:=5mAmph q'#bF5FLFD2_8RI*5HE80-/428E_OFCHO_8IH0RE2+AR5m mpqbh'FL#5F_FDI*2RRH5I8-0E4I2/_FOEH_OCI0H8E+2RR
4;O#FM00NMRb8C0ME_kOl_C#DDRH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2R5b8C04E-2_/8OHEFO8C_CEb02RR+5mAmph q'#bF5FLFD2_IR5*R80CbE2-4/OI_EOFHCC_8b20ER4+R;$
0bFCRkL0_k_#40C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0FjI,RHE80_lMk_DOCD4#-RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0L4k#RF:RkL0_k_#40C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CkRF0k_L#0._$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk.RR:F_k0L.k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#c0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fjc,R*8IH0ME_kOl_C#DD+8dRF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:cRR0Fk_#Lkc$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,UH*I8_0EM_klODCD#R+(8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#U:kRF0k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$LUk#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$LUk#Rb:RN0sH$k_L#0U_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_kn#4_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,4In*HE80_lMk_DOCD4#+6FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4:nRR0Fk_#Lk40n_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bbCRN0sH$k_L#_4n0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#Lk4:nRRsbNH_0$L4k#n$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*d.I0H8Ek_MlC_OD+D#d84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#Rd.:kRF0k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCbHNs0L$_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNbDRN0sH$k_L#Rd.:NRbs$H0_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5b8C0ME_kOl_C#DD-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDHsM_C:oRR8#0_oDFHPO_CFO0sH5I8+0Ed86RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7RQh
o#HMRNDF_k0sRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDF_k0s4CoR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFEROFCF#R0LCIMCCRh7QR8NMR0FkbRk0FAVRD	FORv)q
o#HMRNDs_N8sRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs)7q7)H
#oDMNR8IN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7Wq7#)
HNoMDFRDIN_s8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sd54RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8IN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
o#HMRND)7q7)l_0bRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RbbHCMDHCqR)7
7)#MHoNWDRq)77_b0lR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR7Wq7#)
HNoMDQR7hl_0bRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80bFRHDbCHRMC7
Qh#MHoNWDR l_0bRR:#_08DHFoOR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FbCHbDCHMR
W -C-RML8RD	FORlsNRbHlDCClM00NHRFM#MHoN
D#-L-RCMoHRD#CCRO0sRNlHDlbCMlC0HN0F#MRHNoMDV#
k0MOHRFMo_C0M_kln8c5CEb0:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRNRPD=R:Rb8C0nE/cR;
RRHV5C58bR0ElRF8nRc2>URc2ER0CRM
RPRRN:DR=NRPDRR+4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_knl_cV;
k0MOHRFMo_C0D0CVFsPC_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHL#
CMoH
sRRCs0kMC58bR0ElRF8n;c2
8CMR0oC_VDC0CFPs._d;k
VMHO0FoMRCD0_CFV0P5Cs80CbERR:HCM0o;CsRGlNRH:RMo0CCRs2skC0sHMRMo0CCHsR#N
PsLHNDPCRN:DRR0HMCsoCRR:=jL;
CMoH
HRRV8R5CEb0Rl-RN>GR=2RjRC0EMR
RRNRPD=R:Rb8C0-ERRGlN;R
RCCD#
RRRRDPNRR:=80CbER;
R8CMR;HV
sRRCs0kMN5PD
2;CRM8o_C0D0CVFsPC;k
VMHO0FoMRCM0_kdl_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<c=RUMRN8CR8bR0E>nR42ER0CRM
RRRRPRND:4=R;R
RCRM8H
V;RCRs0MksRDPN;M
C8CRo0k_Ml._d;k
VMHO0FoMRCM0_k4l_nC58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
sPNHDNLCNRPDRR:HCM0oRCs:j=R;C
Lo
HMRVRHRC58bR0E<4=RnMRN8CR8bR0E>2RjRC0EMR
RRPRRN:DR=;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;4n
MOF#M0N0kRMlC_ODnD_cRR:HCM0oRCs:o=RCM0_knl_cC58b20E;F
OMN#0MD0RCFV0P_Csd:.RR0HMCsoCRR:=o_C0D0CVFsPC_5d.80CbE
2;O#FM00NMRlMk_DOCD._dRH:RMo0CC:sR=CRo0k_Ml._d5VDC0CFPs._d2O;
F0M#NRM0D0CVFsPC_R4n:MRH0CCos=R:R0oC_VDC0CFPsC5DVP0FCds_.d,R.
2;O#FM00NMRlMk_DOCDn_4RH:RMo0CC:sR=CRo0k_Mln_45VDC0CFPsn_42
;
0C$bR0Fk_#Lk_b0$Cc_n##RHRsNsN5$RM_klODCD_Rnc8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bCdR.#HN#Rs$sNRk5MlC_ODdD_.FR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$Cn_4##RHRsNsN5$RM_klODCD_R4n8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk_#ncRF:RkL0_k0#_$_bCn;c#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_#d.RF:RkL0_k0#_$_bCd;.#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk_#Lk_#4nRF:RkL0_k0#_$_bC4;n#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$F8VRFRk05bHMk00RFsR0H0-#N#0C2H
#oDMNR0Fk__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-C-RMDNLCV#RF0sRs#H-0CN0#H
#oDMNR0Fk__CMd:.RR8#0_oDFH
O;#MHoNFDRkC0_Mn_4R#:R0D8_FOoH;H
#oDMNR0Is__CM#RR:#_08DHFoOC_POs0F5lMk_DOCDc_nRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-I-RsCH0RNCML#DCRsVFROCNEFRsIVRFRv)qRDOCD##
HNoMDsRI0M_C_Rd.:0R#8F_Do;HO
o#HMRNDI_s0C4M_nRR:#_08DHFoO#;
HNoMDMRH_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-#RkC08RFCRso0H#C7sRQ
hR#MHoNFDRks0_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCs7amz
o#HMRNDs_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDNRI8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDD_FIs8N8sR_#:0R#8F_Do_HOP0COF6s5RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R8N8sHRL0H#RM0bkRR0F)RqvODCD#cR5R0LH#CRsJskHC
82#MHoNDDRFII_Ns88_:#RR8#0_oDFHPO_CFO0sR568MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--Ns88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8-2
-MRC8CR#D0CORlsNRbHlDCClM00NHRFM#MHoN
D#Ns00H0LkC3R\s_NlF#VVCR0\:0R#soHM;L

CMoH
zRRcRd:H5VRs8N8sC_soo2RCsMCNR0C-o-RCsMCNR0CLODF	NRslR
RR-R-RRQVNs88I0H8ERR<OHEFOIC_HE80R#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjjjjjjjjjj&"RR8sN_osC5;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjjjjjj&"RR8IN_osC5;j2
MSC8CRoMNCs0zCRjR;
RzRR4:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjjjjjj&"RR8sN_osC584RF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjjjjj&"RR8IN_osC584RF0IMF2Rj;C
SMo8RCsMCNR0Cz
4;RRRRzR.R:VRHR85N8HsI8R0E=2RdRMoCC0sNCS
SD_FIs8N8s=R<Rj"jjjjjjjjjj&"RR8sN_osC58.RF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjjjjj"RR&I_N8s5Co.FR8IFM0R;j2
MSC8CRoMNCs0zCR.R;
RzRRd:RRRRHV58N8s8IH0=ERRRc2oCCMsCN0
DSSFsI_Ns88RR<="jjjjjjjj"jjRs&RNs8_Cdo5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj&"RR8IN_osC58dRF0IMF2Rj;C
SMo8RCsMCNR0Cz
d;RRRRzRcR:VRHR85N8HsI8R0E=2R6RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjjRj"&NRs8C_soR5c8MFI0jFR2S;
RRRRD_FII8N8s=R<Rj"jjjjjj"jjRI&RNs8_Cco5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR=no2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjj"jjRs&RNs8_C6o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjjjjj"RR&I_N8s5Co6FR8IFM0R;j2
MSC8CRoMNCs0zCR6R;
RzRRn:RRRRHV58N8s8IH0=ERRR(2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjj"jjRs&RNs8_Cno5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj"jjRI&RNs8_Cno5RI8FMR0Fj
2;S8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRNs88I0H8ERR=Uo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjj&"RR8sN_osC58(RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjj"RR&I_N8s5Co(FR8IFM0R;j2
MSC8CRoMNCs0zCR(R;
RzRRU:RRRRHV58N8s8IH0=ERRRg2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjjj&"RR8sN_osC58URF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj"jjRI&RNs8_CUo5RI8FMR0Fj
2;S8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRNs88I0H8ERR=4Rj2oCCMsCN0
RSRRFRDIN_s8R8s<"=Rjjjj"RR&s_N8s5CogFR8IFM0R;j2
DSSFII_Ns88RR<="jjjj&"RR8IN_osC58gRF0IMF2Rj;C
SMo8RCsMCNR0Cz
g;RRRRzR4jRH:RVNR58I8sHE80R4=R4o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jRj"&NRs8C_soj54RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rj"jjRI&RNs8_C4o5jFR8IFM0R;j2
MSC8CRoMNCs0zCR4
j;RRRRzR44RH:RVNR58I8sHE80R4=R.o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC5R448MFI0jFR2S;
SIDF_8IN8<sR=jR"j&"RR8IN_osC5R448MFI0jFR2S;
CRM8oCCMsCN0R4z4;R
RR4Rz.:RRRRHV58N8s8IH0=ERR24dRMoCC0sNCR
SRDRRFsI_Ns88RR<='Rj'&NRs8C_so.54RI8FMR0Fj
2;SFSDIN_I8R8s<'=Rj&'RR8IN_osC5R4.8MFI0jFR2S;
CRM8oCCMsCN0R.z4;R
RR4Rzd:RRRRHV58N8s8IH0>ERR24dRMoCC0sNCR
SRDRRFsI_Ns88RR<=s_N8s5Co48dRF0IMF2Rj;R
SRDRRFII_Ns88RR<=I_N8s5Co48dRF0IMF2Rj;C
SMo8RCsMCNR0Cz;4d
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRcz4RRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<5=R"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj&"RRh7Q2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;S8CMRMoCC0sNC4RzcR;
RzRR4R6R:VRHRF5M0HR8MC_soo2RCsMCN
0CRRRRRRRRRRRRHsM_C<oR="R5jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"RR&72Qh;C
SMo8RCsMCNR0Cz;46
R
RR-R-RRQV5Fs8ks0_CRo2sHCo#s0CR7)_mRzakM#Ho_R)miBp
RRRRnz4RRR:H5VR80Fk_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RmiBp,kRF0C_soR42LHCoMR
RRRRRRRRRRVRHRB5mp=iRR''4R8NMRpmBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRmR7z<aR=kRF0C_so
4;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRRRRRR8CMRMoCC0sNC4RznR;
RzRR4R(R:VRHRF5M0FR8ks0_CRo2oCCMsCN0
RRRRRRRRRRRRz7ma=R<R0Fk_osC4S;
CRM8oCCMsCN0R(z4;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRR4RnsRH:RVsR5Ns88_osC2CRoMNCs0-C
-RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
R--RRRRRRRRRHRRVmR5BRpi=4R''MRN8BRmpCi'P0CM2ER0C-M
-RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
R--RRRRRRRRRCRRMH8RV-;
-RRRRRRRR8CMRFbsO#C#;-
-S8CMRMoCC0sNC4Rzn
s;-R-RR4Rz(:sRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)S;
CRM8oCCMsCN0Rnz4s
;
SR--Q5VRI8N8sC_sos2RC#oH0RCsW7q7)#RkHRMoWB_mpRi
RzRR4RnIRH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8sRCo<W=Rq)7758N8s8IH04E-RI8FMR0Fj
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
MSC8CRoMNCs0zCR4;nI
RRRR(z4IRR:H5VRMRF0I8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRI_N8sRCo<W=Rq)77;C
SMo8RCsMCNR0CzI4(;R

R-RR-GR 0RsNDHFoOFRVskR7NbDRFRs0OCN#
sSzC:oRRFbsO#C#5iBp2CRLo
HMSHRRVBR5p i'ea hR8NMRiBpR'=R4R'20MEC
RSRRh7Q_b0lRR<=7;Qh
RSRR7)q70)_l<bR=qR)7;7)
RSRR7Wq70)_l<bR=qRW7;7)
RSRR_W 0Rlb<W=R S;
RMRC8VRH;C
SMb8RsCFO#
#;
-S-RRQV)8CNR8q8s#C#RW=RsCH0R8q8s#C#,$RLb#N#Rh7QRR0FFbk0kH0RV RWRRH#CLMND
C8SkzlGRR:bOsFC5##W0 _lRb,)7q7)l_0bW,Rq)77_b0l,QR7hl_0bF,Rks0_C
o2SLRRCMoH
RSRRVRHRq5W7_7)0Rlb=qR)7_7)0RlbNRM8W0 _l=bRR''42ER0CSM
SFRRks0_CRo4<7=RQ0h_l
b;SDSC#SC
SFRRks0_CRo4<F=Rks0_CIo5HE80-84RF0IMF2Rj;S
SCRM8H
V;S8CMRFbsO#C#;R
SR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1_
14SUz4RH:RVOR5EOFHCH_I8R0E=2R4RMoCC0sNCR
RRzRS4:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>cR42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR.SzjRR:H5VRNs88I0H8ERR>4Rc2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MR)7q7)l_0b85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24cRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.RzjS;
-Q-RVNR58I8sHE80RR<=4Rc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.4:VRHR85N8HsI8R0E<4=Rco2RCsMCN
0CSSSSF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4z.;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.z.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4Undc7X4RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_d4nU4cX7RR:)Aqv41n_44_1
RSRRRRRRRRRRFRbsl0RN5bR75Qqj=2R>MRH_osC5,[2R7q7)=qR>FRDIN_I858s48dRF0IMF2Rj,QR7A>R=R""j,7Rq7R)A=D>RFsI_Ns885R4d8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5Rj2=F>RkL0_k5#4H2,[2
;
RRRRRRRRRRRRRRRRF_k0s5Co[<2R=kRF0k_L#H45,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
.;RRRRRMSC8CRoMNCs0zCR4
g;RRRRCRM8oCCMsCN0RUz4;RRRRR
RRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_.._1
.SzdRR:H5VROHEFOIC_HE80R.=R2CRoMNCs0RC
RSRRzR.c:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>RdM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRS.:6RRRHV58N8s8IH0>ERR24dRMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM57)q70)_lNb58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMFdR42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCR.
6;SR--Q5VRNs88I0H8E=R<R24dRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRSnz.RH:RVNR58I8sHE80RR<=4Rd2oCCMsCN0
RSRRRRRRRRRRkRF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCR.
n;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRS.:(RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)v4_Ug..X7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)v4_Ug..X7RR:)Aqv41n_.._1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5.[R+48MFI0.FR*,[2R7q7)=qR>FRDIN_I858s48.RF0IMF2Rj,QR7A>R=Rj"j"q,R7A7)RR=>D_FIs8N8s.54RI8FMR0Fj
2,SRSSR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
SSSRRRR7Rmq=F>Rb,CMRA7m5R42=F>RkL0_k5#.H*,.[2+4,mR7A25jRR=>F_k0L.k#5RH,.2*[2R;
RRRRRRRRRRRRRFRRks0_C.o5*R[2<F=RkL0_k5#.H*,.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co.+*[4<2R=kRF0k_L#H.5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCR.
(;RRRRRMSC8CRoMNCs0zCR.
c;RRRRCRM8oCCMsCN0Rdz.;
RR
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11c_cz
S.:URRRHV5FOEH_OCI0H8ERR=co2RCsMCN
0CRRRRSgz.RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4R.2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzRdj:VRHR85N8HsI8R0E>.R42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCR8
RRRRRRRRRRRRRFRRkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR.=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;dj
-S-RRQV58N8s8IH0<ER=.R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSz4RR:H5VRNs88I0H8E=R<R24.RMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';RRRRRRRRRRRRRRRRI_s0CHM52=R<R;W 
RRRRRRRRMSC8CRoMNCs0zCRd
4;SR--tCCMsCN0RC0ERv)qRDOCDN#RM08Rs#H-0CN0#R
RRRRRRzRSd:.RRsVFRH[RMIR5HE80_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqA)vj_cgcnX7RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_cgcnX7RR:)Aqv41n_cc_1
RSRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_so*5c[R+d8MFI0cFR*,[2R7q7)=qR>FRDIN_I858s484RF0IMF2Rj,QR7A>R=Rj"jj,j"R7q7)=AR>FRDIN_s858s484RF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS7Rmq=F>Rb,CMRA7m5Rd2=F>RkL0_k5#cHc,R*d[+27,Rm.A52>R=R0Fk_#Lkc,5Hc+*[.R2,
SSSSA7m5R42=F>RkL0_k5#cH*,c[2+4,mR7A25jRR=>F_k0Lck#5RH,c2*[2R;
RRRRRRRRRRRRRFRRks0_Cco5*R[2<F=RkL0_k5#cH*,c[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[4<2R=kRF0k_L#Hc5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+R.2<F=RkL0_k5#cH*,c[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5c[2+dRR<=F_k0Lck#5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''
;
RRRRRRRRS8CMRMoCC0sNCdRz.R;
RRRRS8CMRMoCC0sNC.RzgR;
RCRRMo8RCsMCNR0Cz;.U
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__1g1Sg
zRdd:VRHRE5OFCHO_8IH0=ERRRg2oCCMsCN0
RRRRdSzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR244RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6zdRH:RVNR58I8sHE80R4>R4o2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4R42=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0R6zd;-
S-VRQR85N8HsI8R0E<4=R4M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSd:nRRRHV58N8s8IH0<ER=4R42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0Rnzd;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS(zdRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv.UjcXRU7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv.UjcXRU7:qR)vnA4__1g1Rg
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[g*+8(RF0IMF*Rg[R2,q)77q>R=RIDF_8IN84s5jFR8IFM0R,j2RA7QRR=>"jjjjjjjjR",q)77A>R=RIDF_8sN84s5jFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBi
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR7Rmq=F>Rb,CMRA7m5R(2=F>RkL0_k5#UH*,U[2+(,mR7A25nRR=>F_k0LUk#5UH,*n[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>kRF0k_L#HU5,[U*+,62RA7m5Rc2=F>RkL0_k5#UH*,U[2+c,mR7A25dRR=>F_k0LUk#5UH,*d[+2
,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.=2R>kRF0k_L#HU5,[U*+,.2RA7m5R42=F>RkL0_k5#UH*,U[2+4,mR7A25jRR=>F_k0LUk#5UH,*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7ujq52>R=R_HMs5Cog+*[UR2,7AQuRR=>",j"Ru7mq>R=RCFbM7,Rm5uAj=2R>NRbs$H0_#LkU,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC5[g*2=R<R0Fk_#LkU,5HU2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+4RR<=F_k0LUk#5UH,*4[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*.[+2=R<R0Fk_#LkU,5HU+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[d<2R=kRF0k_L#HU5,[U*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+Rc2<F=RkL0_k5#UH*,U[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+6RR<=F_k0LUk#5UH,*6[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*n[+2=R<R0Fk_#LkU,5HU+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[(<2R=kRF0k_L#HU5,[U*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+RU2<b=RN0sH$k_L#HU5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRd
(;RRRRRMSC8CRoMNCs0zCRd
c;RRRRCRM8oCCMsCN0Rdzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn4_1U4_1Uz
Sd:URRRHV5FOEH_OCI0H8ERR=4RU2oCCMsCN0
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEM)R5q)77_b0l58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rj2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjzc;-
S-VRQR85N8HsI8R0E<4=RjM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRSc:4RRRHV58N8s8IH0<ER=jR42CRoMNCs0SC
RRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRSRRCRM8oCCMsCN0R4zc;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRS.zcRV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv4cj.X74nRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_.4jcnX47RR:)Aqv41n_41U_4RU
RRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*4U[6+4RI8FMR0F4[U*2q,R7q7)RR=>D_FII8N8sR5g8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858gRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>RpRi,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A6542>R=R0Fk_#Lk4Hn5,*4n[6+427,Rm4A5c=2R>kRF0k_L#54nHn,4*4[+cR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524dRR=>F_k0L4k#n,5H4[n*+24d,mR7A.542>R=R0Fk_#Lk4Hn5,*4n[.+427,Rm4A54=2R>kRF0k_L#54nHn,4*4[+4R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m524jRR=>F_k0L4k#n,5H4[n*+24j,mR7A25gRR=>F_k0L4k#n,5H4[n*+,g2RA7m5RU2=F>RkL0_kn#454H,n+*[UR2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R(2=F>RkL0_kn#454H,n+*[(R2,75mAn=2R>kRF0k_L#54nHn,4*n[+27,Rm6A52>R=R0Fk_#Lk4Hn5,*4n[2+6,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRmcA52>R=R0Fk_#Lk4Hn5,*4n[2+c,mR7A25dRR=>F_k0L4k#n,5H4[n*+,d2RA7m5R.2=F>RkL0_kn#454H,n+*[.R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R42=F>RkL0_kn#454H,n+*[4R2,75mAj=2R>kRF0k_L#54nHn,4*,[2RR
RRRRRRRRRRRRRRRRRRRRRRRRRRQR7u=qR>MRH_osC5*4U[(+4RI8FMR0F4[U*+24n,QR7u=AR>jR"jR",7qmuRR=>FMbC,R
RRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RsbNH_0$L4k#n,5H.+*[4R2,7Amu5Rj2=b>RN0sH$k_L#54nH*,.[;22
RRRRRRRRRRRRRRRR0Fk_osC5*4U[<2R=kRF0k_L#54nHn,4*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+4RR<=F_k0L4k#n,5H4[n*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+.RR<=F_k0L4k#n,5H4[n*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+dRR<=F_k0L4k#n,5H4[n*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+cRR<=F_k0L4k#n,5H4[n*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+6RR<=F_k0L4k#n,5H4[n*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+nRR<=F_k0L4k#n,5H4[n*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+(RR<=F_k0L4k#n,5H4[n*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+URR<=F_k0L4k#n,5H4[n*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[2+gRR<=F_k0L4k#n,5H4[n*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[j+42=R<R0Fk_#Lk4Hn5,*4n[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R42<F=RkL0_kn#454H,n+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[.+42=R<R0Fk_#Lk4Hn5,*4n[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4Rd2<F=RkL0_kn#454H,n+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[c+42=R<R0Fk_#Lk4Hn5,*4n[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R62<F=RkL0_kn#454H,n+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5*4U[n+42=R<RsbNH_0$L4k#n,5H.2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+(<2R=NRbs$H0_#Lk4Hn5,[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRMSC8CRoMNCs0zCRc
.;RRRRRMSC8CRoMNCs0zCRd
g;RRRRCRM8oCCMsCN0RUzd;S

RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAnd_1nd_1nz
SdRUN:VRHRE5OFCHO_8IH0=ERR2dnRMoCC0sNCR
SRzRRdRgN:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80Rg>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
SSSzNcjRH:RVNR58I8sHE80Rg>R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SFSSkC0_M25HRR<='R4'IMECRq5)7_7)05lbNs88I0H8ER-48MFI0gFR2RR=HC2RDR#C';j'
SSSS0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SCSSMo8RCsMCNR0CzNcj;-
S-VRQR85N8HsI8R0E<g=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCS8
ScSz4:NRRRHV58N8s8IH0<ER=2RgRMoCC0sNCS
SSkSF0M_C5RH2<'=R4
';SSSSI_s0CHM52=R<R;W 
SSSCRM8oCCMsCN0R4zcNS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
SSSzNc.RV:RF[sRRRHM58IH0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FAVR)_qv6X4.dR.7:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMS
SS)SAq6v_4d.X.:7RRv)qA_4n1_dn1
dnRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_son5d*d[+4FR8IFM0R*dn[R2,q)77q>R=RIDF_8IN8Us5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5U8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR RRh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,pi
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRq7mRR=>FMbC,mR7A45d2>R=R0Fk_#LkdH.5,*d.[4+d27,RmdA5j=2R>kRF0k_L#5d.H.,d*d[+j
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA.Rg2=F>RkL0_k.#d5dH,.+*[.,g2RA7m52.URR=>F_k0Ldk#.,5Hd[.*+2.U,mR7A(5.2>R=R0Fk_#LkdH.5,*d.[(+.2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm.A5n=2R>kRF0k_L#5d.H.,d*.[+nR2,75mA.R62=F>RkL0_k.#d5dH,.+*[.,62RA7m52.cRR=>F_k0Ldk#.,5Hd[.*+2.c,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7Ad5.2>R=R0Fk_#LkdH.5,*d.[d+.27,Rm.A5.=2R>kRF0k_L#5d.H.,d*.[+.R2,75mA.R42=F>RkL0_k.#d5dH,.+*[.,42
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m52.jRR=>F_k0Ldk#.,5Hd[.*+2.j,mR7Ag542>R=R0Fk_#LkdH.5,*d.[g+427,Rm4A5U=2R>kRF0k_L#5d.H.,d*4[+U
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA4R(2=F>RkL0_k.#d5dH,.+*[4,(2RA7m524nRR=>F_k0Ldk#.,5Hd[.*+24n,mR7A6542>R=R0Fk_#LkdH.5,*d.[6+42R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRm4A5c=2R>kRF0k_L#5d.H.,d*4[+cR2,75mA4Rd2=F>RkL0_k.#d5dH,.+*[4,d2RA7m524.RR=>F_k0Ldk#.,5Hd[.*+24.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7A4542>R=R0Fk_#LkdH.5,*d.[4+427,Rm4A5j=2R>kRF0k_L#5d.H.,d*4[+jR2,75mAg=2R>kRF0k_L#5d.H.,d*g[+2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRmUA52>R=R0Fk_#LkdH.5,*d.[2+U,mR7A25(RR=>F_k0Ldk#.,5Hd[.*+,(2RA7m5Rn2=F>RkL0_k.#d5dH,.+*[n
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR75mA6=2R>kRF0k_L#5d.H.,d*6[+27,RmcA52>R=R0Fk_#LkdH.5,*d.[2+c,mR7A25dRR=>F_k0Ldk#.,5Hd[.*+,d2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRA7m5R.2=F>RkL0_k.#d5dH,.+*[.R2,75mA4=2R>kRF0k_L#5d.H.,d*4[+27,RmjA52>R=R0Fk_#LkdH.5,*d.[
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7qQuRR=>HsM_Cdo5n+*[d86RF0IMFnRd*d[+.R2,7AQuRR=>"jjjjR",7qmuRR=>FMbC,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7udA52>R=RsbNH_0$Ldk#.,5Hc+*[dR2,7Amu5R.2=b>RN0sH$k_L#5d.H*,c[2+.,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRmR7u4A52>R=RsbNH_0$Ldk#.,5Hc+*[4R2,7Amu5Rj2=b>RN0sH$k_L#5d.H*,c[;22
SSSS0Fk_osC5*dn[<2R=kRF0k_L#5d.H.,d*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+4RR<=F_k0Ldk#.,5Hd[.*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+.RR<=F_k0Ldk#.,5Hd[.*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+dRR<=F_k0Ldk#.,5Hd[.*+Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+cRR<=F_k0Ldk#.,5Hd[.*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+6RR<=F_k0Ldk#.,5Hd[.*+R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+nRR<=F_k0Ldk#.,5Hd[.*+Rn2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+(RR<=F_k0Ldk#.,5Hd[.*+R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+URR<=F_k0Ldk#.,5Hd[.*+RU2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[2+gRR<=F_k0Ldk#.,5Hd[.*+Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+42=R<R0Fk_#LkdH.5,*d.[j+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R42<F=RkL0_k.#d5dH,.+*[4R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+42=R<R0Fk_#LkdH.5,*d.[.+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4Rd2<F=RkL0_k.#d5dH,.+*[4Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+42=R<R0Fk_#LkdH.5,*d.[c+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R62<F=RkL0_k.#d5dH,.+*[4R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[n+42=R<R0Fk_#LkdH.5,*d.[n+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4R(2<F=RkL0_k.#d5dH,.+*[4R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[U+42=R<R0Fk_#LkdH.5,*d.[U+42ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[4Rg2<F=RkL0_k.#d5dH,.+*[4Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+.2=R<R0Fk_#LkdH.5,*d.[j+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R42<F=RkL0_k.#d5dH,.+*[.R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+.2=R<R0Fk_#LkdH.5,*d.[.+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.Rd2<F=RkL0_k.#d5dH,.+*[.Rd2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+.2=R<R0Fk_#LkdH.5,*d.[c+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R62<F=RkL0_k.#d5dH,.+*[.R62IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[n+.2=R<R0Fk_#LkdH.5,*d.[n+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.R(2<F=RkL0_k.#d5dH,.+*[.R(2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[U+.2=R<R0Fk_#LkdH.5,*d.[U+.2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[.Rg2<F=RkL0_k.#d5dH,.+*[.Rg2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[j+d2=R<R0Fk_#LkdH.5,*d.[j+d2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[dR42<F=RkL0_k.#d5dH,.+*[dR42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[.+d2=R<RsbNH_0$Ldk#.,5Hc2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+d<2R=NRbs$H0_#LkdH.5,[c*+R42IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[c+d2=R<RsbNH_0$Ldk#.,5Hc+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2d6RR<=bHNs0L$_k.#d5cH,*d[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SMSC8CRoMNCs0zCRc;.N
CSSMo8RCsMCNR0CzNdg;C
SMo8RCsMCNR0CzNdU;R
RCRM8oCCMsCN0Rdzc;R

RczcRH:RVMR5Fs0RNs88_osC2CRoMNCs0-CR-CRoMNCs0#CRCODC0NRslR
RR-R-RRQVNs88I0H8ERR<6#RN#MHoR''jRR0Fk#MkCL8RH
0#RRRRzRjR:VRHR85N8HsI8R0E=2R4RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jj"jjRs&RNs8_C#o_5;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjjRj"&NRI8C_so5_#j
2;RRRRCRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j"jjRs&RNs8_C#o_584RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jjRj"&NRI8C_so5_#4FR8IFM0R;j2
RRRR8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<"=Rj"jjRs&RNs8_C#o_58.RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<Rj"jj&"RR8IN_osC_.#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"j&"RR8sN_osC_d#5RI8FMR0Fj
2;RRRRRRRRD_FII8N8sR_#<"=RjRj"&NRI8C_so5_#dFR8IFM0R;j2
RRRR8CMRMoCC0sNCdRz;z
ScRS:H5VRNs88I0H8ERR=6o2RCsMCN
0CSFSDIN_s8_8s#=R<R''jRs&RNs8_C#o_58cRF0IMF2Rj;S
SD_FII8N8sR_#<'=Rj&'RR8IN_osC_c#5RI8FMR0Fj
2;S8CMRMoCC0sNCcRz;R
RR6RzRRR:H5VRNs88I0H8ERR>6o2RCsMCN
0CRRRRRRRRD_FIs8N8sR_#<s=RNs8_C#o_586RF0IMF2Rj;R
RRRRRRFRDIN_I8_8s#=R<R8IN_osC_6#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z6
R
RR-R-RRQV5M8H_osC2CRso0H#C7sRQkhR#oHMRiBp
RRRRRznRH:RV8R5HsM_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5Bi7,RQRh2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRHsM_C#o_RR<=7;Qh
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRnR;
RzRR(:RRRRHV50MFRM8H_osC2CRoMNCs0RC
RRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRCRM8oCCMsCN0R;z(
R
RR-R-RRQV5k8F0C_sos2RC#oH0RCs7amzRHk#MmoRB
piRRRRzRUR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s_Co#L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRRz7ma=R<R0Fk_osC_
#;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCURz;R
RRgRzRRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C#o_;R
RRMRC8CRoMNCs0zCRg
;
RRRR-Q-RVNR58_8ss2CoRosCHC#0s7Rq7k)R#oHMRiBp
RRRRjz4RRR:H5VRs8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qR)727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osC_<#R=qR)757)Ns88I0H8ER-48MFI0jFR2R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0Rjz4;R
RR4Rz4RR:H5VRMRF0s8N8sC_soo2RCsMCN
0CRRRRRRRRRRRRs_N8s_Co#=R<R7)q7
);RRRRCRM8oCCMsCN0R4z4;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4.RH:RVIR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7Wq7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRI_N8s_Co#=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4.
RRRRdz4RH:RVMR5FI0RNs88_osC2CRoMNCs0RC
RRRRRRRRRIRRNs8_C#o_RR<=W7q7)R;
RCRRMo8RCsMCNR0Cz;4d
RRRRRRRRR
RR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoH
RRRRcz4RV:RFHsRRRHM5lMk_DOCDc_nR4-R2FR8IFM0RojRCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRR6z4RH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M5_#H<2R=4R''ERIC5MRs_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RWRCIEMIR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4
6;RRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR4n:VRHR85N8HsI8R0E<n=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M5_#H<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M5_#H<2R= RW;R
RRRRRRMRC8CRoMNCs0zCR4
n;RRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR(z4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRnc:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNC*5HnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05+5H4n2*c8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRnc:)RXqcvnXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RRq6=D>RFII_Ns88_6#52
,RSSSSSRSR7qu)j>R=RIDF_8sN8#s_5,j2R)7uq=4R>FRDIN_s8_8s#254,uR7)Rq.=D>RFsI_Ns88_.#52S,
SSSSS7RRud)qRR=>D_FIs8N8s5_#dR2,7qu)c>R=RIDF_8sN8#s_5,c2R)7uq=6R>FRDIN_s8_8s#256,SR
SSSSSWRR >R=R0Is__CM#25H,BRWp=iR>pRBi7,Ru=mR>kRF0k_L#c_n#,5H[;22
RRRRRRRRRRRRRRRR0Fk_osC_[#52=R<R0Fk_#Lk_#nc5[H,2ERIC5MRF_k0C#M_5RH2=4R''C2RDR#C';Z'
RRRRRRRR8CMRMoCC0sNC4Rz(R;
RRRRCRM8oCCMsCN0Rcz4;RRRRRRRRRRRRR
RRRRR
RRRRR--tCCMsCN0RdNR.FRIs88RCRCb)RqvODCDRRHVNsbbFHbsNR0CRRRRRRRRRRRRRRR
RzRR4:URRRHV5lMk_DOCD._dR4=R2CRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R(RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzN4gRH:RVNR58I8sHE80Rn>R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rgz4NR;
RRRRRzRR4RgL:VRHR85N8HsI8R0E=RRnNRM8M_klODCD_Rnc=2RjRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5N5s8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzL4g;RRRRR--Q5VRNs88I0H8E=R<RR62MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRjz.RH:RVNR58I8sHE80RR<=6o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CdM_.=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_Rd.<W=R R;
RRRRRCRRMo8RCsMCNR0Cz;.j
RRRRR--tCCMsCN0RC0ERv)qRDOCDMRN8sR0H0-#N
0CRRRRRRRRzR.4:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qd:.RRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5lMk_DOCDc_n*2ncR"&RW&"RR0HMCsoC'NHlo[C52RR&"R "&MRH0CCosl'HN5oCo_C0C_M880CbEk5MlC_ODnD_cc*nRd+R.8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vRd.:)RXq.vdXR47
RRRRRRRRRRRRRRRRsbF0NRlb7R5RR=>HsM_C#o_5,[2RRqj=D>RFII_Ns88_j#52q,R4>R=RIDF_8IN8#s_5,42RRq.=D>RFII_Ns88_.#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRRqd=D>RFII_Ns88_d#52q,Rc>R=RIDF_8IN8#s_5,c2RS
SSSSSRuR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d,uR7)Rqc=D>RFsI_Ns88_c#52
,RSSSSSRSRW= R>sRI0M_C_,d.RpWBi>R=RiBp,uR7m>R=R0Fk_#Lk_#d.5lMk_DOCD._d,2[2;R
RRRRRRRRRRRRRRkRF0C_so5_#[<2R=kRF0k_L#._d#k5MlC_ODdD_.2,[RCIEMFR5kC0_M._dR'=R4R'2CCD#R''Z;R
RRRRRRCRRMo8RCsMCNR0Cz;.4
RRRRMRC8CRoMNCs0zCR4RU;RRRRRRRRRR

R-RR-CRtMNCs0NCRRR4nI8FsRC8CbqR)vCRODHDRVbRNbbsFs0HNCRRRRRRRRRRRRRRR
RRRR.z.RH:RVMR5kOl_C_DD4=nRRR42oCCMsCN0
RRRRR--Q5VRNs88I0H8ERR>6M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR.Rzd:NRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd=.RRR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858sN_osC_6#52RR='24'R8NMRN5s8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CM4<nR= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=R4R'2NRM858IN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.NR;
RRRRRzRR.RdL:VRHR85N8HsI8R0E>RRnNRM8M_klODCD_Rd./4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8sR5Ns8_C#o_5R62=jR''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5I8C_so5_#6=2RR''j2MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dL
RRRRRRRRdz.ORR:H5VRNs88I0H8ERR=nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzO.d;R
RRRRRR.Rzd:8RRRHV58N8s8IH0=ERRN6RMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fc=2RRlMk_DOCD._d2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.RzdR8;R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR.:cRRRHV58N8s8IH0<ER=2RcRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<R;W 
RRRRRRRR8CMRMoCC0sNC.RzcR;
R-RR-CRtMNCs00CRE)CRqOvRCRDDNRM80-sH#00NCR
RRRRRR.Rz6RR:VRFs[MRHRH5I8R0E-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)Rzqnv4RD:RNDLCRRH#"a17"RR&HCM0o'CsHolNCH5I820ER"&R7&"RR0HMCsoC'NHloMC5kOl_C_DDnnc*cRR+M_klODCD_*d.dR.2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+kRMlC_ODdD_..*dR4+Rn8,RCEb02&2RR""XRH&RMo0CCHs'lCNo54[+2R;
RRRRRRRRRLRRCMoH
RRRRRRRRRRRRqz)vR4n:qR)vX4n4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,uR7)Rqj=D>RFsI_Ns88_j#527,Ru4)qRR=>D_FIs8N8s5_#4R2,7qu).>R=RIDF_8sN8#s_5,.2
SSSSRSSR)7uq=dR>FRDIN_s8_8s#25d, RWRR=>I_s0C4M_nW,RBRpi=B>RpRi,7Rum=F>RkL0_k4#_nM#5kOl_C_DD4[n,2
2;RRRRRRRRRRRRRRRRF_k0s_Co#25[RR<=F_k0L_k#45n#M_klODCD_,4n[I2RERCM50Fk__CM4=nRR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R6z.;R
RRMRC8CRoMNCs0zCR.R.;R
RRRMRC8CRoMNCs0zCRc
c;CRM8NEsOHO0C0CksRFLDOs	_N
l;
ONsECH0Os0kCFRM__sIOOEC	VRFRv)q_W)_R
H#ObFlFMMC0)RXq.vdXR47RFRbs50R
RRRRRRRRm7uR:RRR0FkR8#0_FkDo;HORRRRRRRR
RRRRRRRRm1uR:RRR0FkR8#0_FkDo;HO
R
RRRRRRjRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRq4R:RRRRHM#_08koDFH
O;RRRRRRRRqR.RRRR:H#MR0k8_DHFoOR;
RRRRRqRRdRRRRH:RM0R#8D_kFOoH;R
RRRRRRcRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRR7RR:RRRRHM#_08koDFH
O;RRRRRRRR7qu)jRR:H#MR0k8_DHFoOR;
RRRRR7RRu4)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rq.:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:dRRRHM#_08koDFH
O;RRRRRRRR7qu)cRR:H#MR0k8_DHFoOR;
RRRRRWRRBRpiRH:RM0R#8D_kFOoH;RRRRRRRRR
RRRRRR RWRRRR:MRHR8#0_FkDo
HORRRRR2RR;
RRCRM8ObFlFMMC0O;
FFlbM0CMRqX)vXnc4R7RRsbF0
R5RRRRRRRR7RumRRR:FRk0#_08koDFHRO;RRRRR
RRRRRRRRRR1RumRRR:FRk0#_08koDFH
O;
RRRRRRRRRqjR:RRRRHM#_08koDFH
O;RRRRRRRRqR4RRRR:H#MR0k8_DHFoOR;
RRRRRqRR.RRRRH:RM0R#8D_kFOoH;R
RRRRRRdRqRRRR:MRHR8#0_FkDo;HO
RRRRRRRRRqcR:RRRRHM#_08koDFH
O;RRRRRRRRqR6RRRR:H#MR0k8_DHFoOR;
RRRRR7RRRRRRRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqj:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:4RRRHM#_08koDFH
O;RRRRRRRR7qu).RR:H#MR0k8_DHFoOR;
RRRRR7RRud)qRH:RM0R#8D_kFOoH;R
RRRRRRuR7)Rqc:MRHR8#0_FkDo;HO
RRRRRRRR)7uq:6RRRHM#_08koDFH
O;RRRRRRRRWiBpRRR:H#MR0k8_DHFoOR;RRRRRRRR
RRRRRWRR RRRRH:RM0R#8D_kFOoH
RRRRRRR2R;R
8CMRlOFbCFMM
0;VOkM0MHFRMVkOM_HHL05RL:RFCFDNRM2skC0s#MR0MsHo#RH
oLCHRM
RRHV5RL20MEC
RRRR0sCk5sM"RhFs8CN/HIs0OCRFDMVHRO0OOEC	13RHDlkNF0HMHRl#0lNObERFH##LRDC!2!";R
RCCD#
RRRR0sCk5sM"kBFDM8RFH0RlCbDl0CMRFADO)	RqRv3Q0#REsCRCRN8Ns88CR##sHCo#s0CCk8R#oHMRC0ERl#NCDROFRO	N0#RE)CRq"v?2R;
R8CMR;HV
8CMRMVkOM_HH
0;VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEN;
0H0sLCk0RMoCC0sNFss_CsbF0RR:#H0sM
o;Ns00H0LkCCRoMNCs0_FssFCbsF0RVFRM__sIOOEC	RR:NEsOHO0C0CksRRH#VOkM_HHM0N5s8_8ss2Co;-
-RoLCHLMRD	FORlsNRbHlDCClM00NHRFM#MHoN
D#0C$bR0HM_sNsNH$R#sRNsRN$50jRF2R6RRFVHCM0o;Cs
MOF#M0N0HRI8_0ENNss$RR:H_M0NNss$=R:R,54RR.,cg,R,UR4,nRd2O;
F0M#NRM080CbEs_NsRN$:MRH0s_NsRN$:5=R4UndcU,R4,g.Rgcjn.,Rj,cUR.4jc6,R4;.2
MOF#M0N0HR8PRd.:MRH0CCos=R:RH5I8-0E4d2/nO;
F0M#NRM084HPnRR:HCM0oRCs:5=RI0H8E2-4/;4U
MOF#M0N0HR8P:URR0HMCsoCRR:=58IH04E-2;/g
MOF#M0N0HR8P:cRR0HMCsoCRR:=58IH04E-2;/c
MOF#M0N0HR8P:.RR0HMCsoCRR:=58IH04E-2;/.
MOF#M0N0HR8P:4RR0HMCsoCRR:=58IH04E-2;/4
F
OMN#0ML0RF4FDRL:RFCFDN:MR=8R5HRP4>2Rj;F
OMN#0ML0RF.FDRL:RFCFDN:MR=8R5HRP.>2Rj;F
OMN#0ML0RFcFDRL:RFCFDN:MR=8R5HRPc>2Rj;F
OMN#0ML0RFUFDRL:RFCFDN:MR=8R5HRPU>2Rj;F
OMN#0ML0RF4FDnRR:LDFFCRNM:5=R84HPnRR>j
2;O#FM00NMRFLFDRd.:FRLFNDCM=R:RH58PRd.>2Rj;O

F0M#NRM084HPncdURH:RMo0CC:sR=8R5CEb0-/424UndcO;
F0M#NRM08UHP4Rg.:MRH0CCos=R:RC58b-0E4U2/4;g.
MOF#M0N0HR8PgcjnRR:HCM0oRCs:5=R80CbE2-4/gcjnO;
F0M#NRM08.HPjRcU:MRH0CCos=R:RC58b-0E4.2/j;cU
MOF#M0N0HR8P.4jcRR:HCM0oRCs:5=R80CbE2-4/.4jcO;
F0M#NRM086HP4:.RR0HMCsoCRR:=5b8C04E-24/6.
;
O#FM00NMRFLFD.64RL:RFCFDN:MR=8R5H4P6.RR>j
2;O#FM00NMRFLFD.4jcRR:LDFFCRNM:5=R84HPjR.c>2Rj;F
OMN#0ML0RF.FDjRcU:FRLFNDCM=R:RH58Pc.jURR>j
2;O#FM00NMRFLFDgcjnRR:LDFFCRNM:5=R8cHPjRgn>2Rj;F
OMN#0ML0RFUFD4Rg.:FRLFNDCM=R:RH58PgU4.RR>j
2;O#FM00NMRFLFDd4nU:cRRFLFDMCNRR:=5P8H4UndcRR>j
2;
MOF#M0N0kR#lH_I8R0E:MRH0CCos=R:RmAmph q'#bF5FLFDR42+mRAmqp hF'b#F5LF2D.RA+Rm mpqbh'FL#5FcFD2RR+Apmm 'qhb5F#LDFFU+2RRmAmph q'#bF5FLFD24n;F
OMN#0M#0Rk8l_CEb0RH:RMo0CC:sR=RR6-AR5m mpqbh'FL#5F6FD4R.2+mRAmqp hF'b#F5LFjD4.Rc2+mRAmqp hF'b#F5LFjD.cRU2+mRAmqp hF'b#F5LFjDcgRn2+mRAmqp hF'b#F5LF4DUg2.2;O

F0M#NRM0IE_OFCHO_8IH0:ERR0HMCsoCRR:=I0H8Es_Ns5N$#_klI0H8E
2;O#FM00NMROI_EOFHCC_8bR0E:MRH0CCos=R:Rb8C0NE_s$sN5l#k_8IH0;E2
MOF#M0N0_R8OHEFOIC_HE80RH:RMo0CC:sR=HRI8_0ENNss$k5#lC_8b20E;F
OMN#0M80R_FOEH_OC80CbERR:HCM0oRCs:8=RCEb0_sNsN#$5k8l_CEb02
;
O#FM00NMRII_HE80_lMk_DOCD:#RR0HMCsoCRR:=58IH04E-2_/IOHEFOIC_HE80R4+R;F
OMN#0MI0R_b8C0ME_kOl_C#DDRH:RMo0CC:sR=8R5CEb0-/42IE_OFCHO_b8C0+ERR
4;
MOF#M0N0_R8I0H8Ek_MlC_ODRD#:MRH0CCos=R:RH5I8-0E482/_FOEH_OCI0H8ERR+4O;
F0M#NRM08C_8b_0EM_klODCD#RR:HCM0oRCs:5=R80CbE2-4/O8_EOFHCC_8bR0E+;R4
F
OMN#0MI0R_x#HCRR:HCM0oRCs:I=R_8IH0ME_kOl_C#DDRI*R_b8C0ME_kOl_C#DD;F
OMN#0M80R_x#HCRR:HCM0oRCs:8=R_8IH0ME_kOl_C#DDR8*R_b8C0ME_kOl_C#DD;O

F0M#NRM0LDFF_:8RRFLFDMCNRR:=5#8_HRxC-_RI#CHxRR<=j
2;O#FM00NMRFLFDR_I:FRLFNDCM=R:R0MF5FLFD2_8;O

F0M#NRM0OHEFOIC_HE80RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFOIC_HE802O;
F0M#NRM0OHEFO8C_CEb0RH:RMo0CC:sR=AR5m mpqbh'FL#5F_FD8*2RRO8_EOFHCC_8b20ER5+RApmm 'qhb5F#LDFF_RI2*_RIOHEFO8C_CEb02O;
F0M#NRM0I0H8Ek_MlC_ODRD#:MRH0CCos=R:Rm5Amqp hF'b#F5LF8D_25R*I0H8E2-4/O8_EOFHCH_I820ER5+RApmm 'qhb5F#LDFF_RI2*IR5HE80-/42IE_OFCHO_8IH0RE2+;R4
MOF#M0N0CR8b_0EM_klODCD#RR:HCM0oRCs:5=RApmm 'qhb5F#LDFF_R82*C58b-0E482/_FOEH_OC80CbE+2RRm5Amqp hF'b#F5LFID_2RR*5b8C04E-2_/IOHEFO8C_CEb02RR+40;
$RbCF_k0L4k#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,I0H8Ek_MlC_OD-D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lk4RR:F_k0L4k#_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k_#.0C$bRRH#NNss$8R5CEb0_lMk_DOCD4#-RI8FMR0Fj.,R*8IH0ME_kOl_C#DD+84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#:.RR0Fk_#Lk.$_0bRC;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0Lck#_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,cH*I8_0EM_klODCD#R+d8MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kR#c:kRF0k_L#0c_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bR0Fk_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIU*HE80_lMk_DOCD(#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDF_k0LUk#RF:RkL0_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#LkU$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR8IH0ME_kOl_C#DD-84RF0IMF2RjRRFV#_08DHFoO#;
HNoMDNRbs$H0_#LkURR:bHNs0L$_k_#U0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RV_Rs80FkRM5HbRk000FRs#H-0CN0#02
$RbCF_k0L4k#n$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjR*4nI0H8Ek_MlC_OD+D#486RF0IMF2RjRRFV#_08DHFoO#;
HNoMDkRF0k_L#R4n:kRF0k_L#_4n0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
b0$CNRbs$H0_#Lk40n_$RbCHN#Rs$sNRC58b_0EM_klODCD#R-48MFI0jFR,*R.I0H8Ek_MlC_OD+D#4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNRsbNH_0$L4k#nRR:bHNs0L$_kn#4_b0$CR;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFR8s_FRk05bHMk00RFsR0H0-#N#0C2$
0bFCRkL0_k.#d_b0$C#RHRsNsN5$R80CbEk_MlC_OD-D#4FR8IFM0RRj,dI.*HE80_lMk_DOCDd#+4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#Lkd:.RR0Fk_#Lkd0._$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-.-R7sRNsRN$FsVR_k8F0HR5M0bkRR0F0-sH#00NC
#20C$bRsbNH_0$Ldk#.$_0bHCR#sRNsRN$5b8C0ME_kOl_C#DD-84RF0IMF,RjRIc*HE80_lMk_DOCDd#+RI8FMR0FjF2RV0R#8F_Do;HO
o#HMRNDbHNs0L$_k.#dRb:RN0sH$k_L#_d.0C$b;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--.N7Rs$sNRRFVsF_8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRCNCLD#FRVssR0H0-#N#0C
o#HMRNDI_s0C:MRR8#0_oDFHPO_CFO0sC58b_0EM_klODCD#R-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRIHR0CCLMNDRC#VRFsCENORIsFRRFV)RqvODCD#H
#oDMNR_HMsRCo:0R#8F_Do_HOP0COFIs5HE80+Rd68MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8E6+dRI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRz7maH
#oDMNR0Fk_osC4RR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80OFRE#FFCCRL0CICMQR7hMRN8kRF00bkRRFVAODF	qR)vH
#oDMNR8sN_osCR#:R0D8_FOoH_OPC05FsNs88I0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0sqRW7
7)#MHoNDDRFsI_Ns88R#:R0D8_FOoH_OPC05Fs48dRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RNs88R0LH#MRHbRk00)FRqOvRC#DDRR5cL#H0RJsCkCHs8#2
HNoMDFRDIN_I8R8s:0R#8F_Do_HOP0COF4s5dFR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRNs_8_8ssRCo:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;-
-R8CMRFLDOs	RNHlRlCbDl0CMNF0HMHR#oDMN#-
-RoLCH#MRCODC0NRsllRHblDCCNM00MHFRo#HM#ND
MVkOF0HMCRo0k_Mlc_n5b8C0RE:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RPRND:8=RCEb0/;nc
HRRV5R580CbEFRl8cRn2RR>cRU20MEC
RRRRDPNRR:=PRND+;R4
CRRMH8RVR;
R0sCkRsMP;ND
8CMR0oC_lMk_;nc
MVkOF0HMCRo0C_DVP0FCds_.C58bR0E:MRH0CCoss2RCs0kMMRH0CCos#RH
oLCHRM
R0sCk5sM80CbEFRl8cRn2C;
Mo8RCD0_CFV0P_Csd
.;VOkM0MHFR0oC_VDC0CFPsC58bR0E:MRH0CCosl;RN:GRR0HMCsoC2CRs0MksR0HMCsoCR
H#PHNsNCLDRDPNRH:RMo0CC:sR=;Rj
oLCHRM
RRHV5b8C0-ERRGlNRR>=j02RE
CMRRRRPRND:8=RCEb0Rl-RN
G;RDRC#RC
RPRRN:DR=CR8b;0E
CRRMH8RVR;
R0sCk5sMP2ND;M
C8CRo0C_DVP0FC
s;VOkM0MHFR0oC_lMk_5d.80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RRcUNRM880CbERR>4Rn20MEC
RRRRNRPD=R:R
4;RMRC8VRH;R
RskC0sPMRN
D;CRM8o_C0M_kld
.;VOkM0MHFR0oC_lMk_54n80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCPRND:MRH0CCos=R:R
j;LHCoMR
RH5VR80CbE=R<RR4nNRM880CbERR>j02RE
CMRRRRRDPNRR:=4R;
R8CMR;HV
sRRCs0kMNRPDC;
Mo8RCM0_k4l_nO;
F0M#NRM0M_klODCD_Rnc:MRH0CCos=R:R0oC_lMk_5nc80CbE
2;O#FM00NMRVDC0CFPs._dRH:RMo0CC:sR=CRo0C_DVP0FCds_.C58b20E;F
OMN#0MM0RkOl_C_DDd:.RR0HMCsoCRR:=o_C0M_kldD.5CFV0P_Csd;.2
MOF#M0N0CRDVP0FC4s_nRR:HCM0oRCs:o=RCD0_CFV0P5CsD0CVFsPC_,d.R2d.;F
OMN#0MM0RkOl_C_DD4:nRR0HMCsoCRR:=o_C0M_kl4Dn5CFV0P_Cs4;n2
$
0bFCRkL0_k0#_$_bCnRc#HN#Rs$sNRk5MlC_ODnD_cFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;0C$bR0Fk_#Lk_b0$C._d##RHRsNsN5$RM_klODCD_Rd.8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;$
0bFCRkL0_k0#_$_bC4Rn#HN#Rs$sNRk5MlC_OD4D_nFR8IFM0RRj,I0H8ER-48MFI0jFR2VRFR8#0_oDFH
O;#MHoNFDRkL0_kn#_c:#RR0Fk_#Lk_b0$Cc_n#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_kd#_.:#RR0Fk_#Lk_b0$C._d#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkL0_k4#_n:#RR0Fk_#Lk_b0$Cn_4#R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RR.7NNss$VRFRk8F0HR5M0bkRR0F0-sH#00NC
#2#MHoNFDRkC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNFDRkC0_M._dR#:R0D8_FOoH;H
#oDMNR0Fk__CM4:nRR8#0_oDFH
O;#MHoNIDRsC0_MR_#:0R#8F_Do_HOP0COFMs5kOl_C_DDn8cRF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RHIs0CCRMDNLCV#RFCsRNROEsRFIF)VRqOvRC#DD
o#HMRNDI_s0CdM_.RR:#_08DHFoO#;
HNoMDsRI0M_C_R4n:0R#8F_Do;HO
o#HMRNDHsM_C#o_R#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osC_:#RR8#0_oDFHPO_CFO0sH5I8-0E4FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0smR7z#a
HNoMDNRs8C_soR_#:0R#8F_Do_HOP0COFNs58I8sHE80-84RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-k-R#RC80sFRC#oH0RCsq)77
o#HMRNDI_N8s_Co#RR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCk#8FR0RosCHC#0s7Rq7#)
HNoMDFRDIN_s8_8s#RR:#_08DHFoOC_POs0F586RF0IMF2Rj;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-N-R8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8#s_R#:R0D8_FOoH_OPC05Fs6FR8IFM0R;j2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-8RN8LsRHR0#HkMb0FR0Rv)qRDOCD5#RcHRL0s#RCHJks2C8
R--CRM8#CCDOs0RNHlRlCbDl0CMNF0HMHR#oDMN#0
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCHRM
Rdzc:VRHRN5s8_8ss2CoRMoCC0sNC-R-RMoCC0sNCDRLFRO	s
NlRRRR-Q-RV8RN8HsI8R0E<EROFCHO_8IH0NER#o#HMjR''FR0RkkM#RC8L#H0
RRRRRzjRH:RVNR58I8sHE80R4=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjjjjjj"jjRs&RNs8_Cjo52S;
RRRRD_FII8N8s=R<Rj"jjjjjjjjjj"jjRI&RNs8_Cjo52S;
CRM8oCCMsCN0R;zj
RRRRRz4RH:RVNR58I8sHE80R.=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj"jjRs&RNs8_C4o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjj"jjRI&RNs8_C4o5RI8FMR0Fj
2;S8CMRMoCC0sNC4Rz;R
RR.RzRRR:H5VRNs88I0H8ERR=do2RCsMCN
0CSFSDIN_s8R8s<"=Rjjjjjjjjj"jjRs&RNs8_C.o5RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=jR"jjjjjjjjjRj"&NRI8C_soR5.8MFI0jFR2S;
CRM8oCCMsCN0R;z.
RRRRRzdRH:RVNR58I8sHE80Rc=R2CRoMNCs0SC
SIDF_8sN8<sR=jR"jjjjjjjjj&"RR8sN_osC58dRF0IMF2Rj;R
SRDRRFII_Ns88RR<="jjjjjjjj"jjRI&RNs8_Cdo5RI8FMR0Fj
2;S8CMRMoCC0sNCdRz;R
RRcRzRRR:H5VRNs88I0H8ERR=6o2RCsMCN
0CSRRRRIDF_8sN8<sR=jR"jjjjjjjj"RR&s_N8s5CocFR8IFM0R;j2
RSRRFRDIN_I8R8s<"=Rjjjjjjjjj&"RR8IN_osC58cRF0IMF2Rj;C
SMo8RCsMCNR0Cz
c;RRRRzR6R:VRHR85N8HsI8R0E=2RnRMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjjjjjj&"RR8sN_osC586RF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjjRj"&NRI8C_soR568MFI0jFR2S;
CRM8oCCMsCN0R;z6
RRRRRznRH:RVNR58I8sHE80R(=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjjjjj&"RR8sN_osC58nRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jjjjjj&"RR8IN_osC58nRF0IMF2Rj;C
SMo8RCsMCNR0Cz
n;RRRRzR(R:VRHR85N8HsI8R0E=2RURMoCC0sNCR
SRDRRFsI_Ns88RR<="jjjj"jjRs&RNs8_C(o5RI8FMR0Fj
2;SFSDIN_I8R8s<"=RjjjjjRj"&NRI8C_soR5(8MFI0jFR2S;
CRM8oCCMsCN0R;z(
RRRRRzURH:RVNR58I8sHE80Rg=R2CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jj"jjRs&RNs8_CUo5RI8FMR0Fj
2;SFSDIN_I8R8s<"=Rjjjjj&"RR8IN_osC58URF0IMF2Rj;C
SMo8RCsMCNR0Cz
U;RRRRzRgR:VRHR85N8HsI8R0E=jR42CRoMNCs0SC
RRRRD_FIs8N8s=R<Rj"jjRj"&NRs8C_soR5g8MFI0jFR2S;
SIDF_8IN8<sR=jR"j"jjRI&RNs8_Cgo5RI8FMR0Fj
2;S8CMRMoCC0sNCgRz;R
RR4Rzj:RRRRHV58N8s8IH0=ERR244RMoCC0sNCR
SRDRRFsI_Ns88RR<="jjj"RR&s_N8s5Co48jRF0IMF2Rj;S
SD_FII8N8s=R<Rj"jj&"RR8IN_osC5R4j8MFI0jFR2S;
CRM8oCCMsCN0Rjz4;R
RR4Rz4:RRRRHV58N8s8IH0=ERR24.RMoCC0sNCR
SRDRRFsI_Ns88RR<=""jjRs&RNs8_C4o54FR8IFM0R;j2
DSSFII_Ns88RR<=""jjRI&RNs8_C4o54FR8IFM0R;j2
MSC8CRoMNCs0zCR4
4;RRRRzR4.RH:RVNR58I8sHE80R4=Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=jR''RR&s_N8s5Co48.RF0IMF2Rj;S
SD_FII8N8s=R<R''jRI&RNs8_C4o5.FR8IFM0R;j2
MSC8CRoMNCs0zCR4
.;RRRRzR4dRH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSRRRRIDF_8sN8<sR=NRs8C_sod54RI8FMR0Fj
2;SRRRRIDF_8IN8<sR=NRI8C_sod54RI8FMR0Fj
2;S8CMRMoCC0sNC4Rzd
;
RRRR-Q-RV8R5HsM_CRo2sHCo#s0CRh7QRHk#MBoRpRi
RzRR4RcR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_so=R<Rj5"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jjR7&RQ;h2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;C
SMo8RCsMCNR0Cz;4c
RRRR6z4RRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=5j"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjRj"&QR7h
2;S8CMRMoCC0sNC4Rz6
;
RRRR-Q-RVsR580Fk_osC2CRso0H#C)sR_z7ma#RkHRMo)B_mpRi
RzRR4RnR:VRHRF58ks0_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,F_k0s4Co2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s4Co;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RRRRRCRRMo8RCsMCNR0Cz;4n
RRRR(z4RRR:H5VRMRF080Fk_osC2CRoMNCs0RC
RRRRRRRRR7RRmRza<F=Rks0_C;o4
MSC8CRoMNCs0zCR4
(;
RRRRR--Q5VRs8N8sC_sos2RC#oH0RCs)7q7)#RkHRMomiBp
RRRRnz4s:RRRRHV58sN8ss_CRo2oCCMsCN0
R--RRRRRbRRsCFO#5#RmiBp,qR)727)RoLCH-M
-RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
R--RRRRRRRRRRRRRsRRNs8_C<oR=qR)757)Ns88I0H8ER-48MFI0jFR2-;
-RRRRRRRRRRRR8CMR;HV
R--RRRRRCRRMb8RsCFO#
#;-C-SMo8RCsMCNR0Czs4n;-
-RRRRzs4(RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C<oR=qR)7;7)
MSC8CRoMNCs0zCR4;ns
-
S-VRQRN5I8_8ss2CoRosCHC#0sqRW7R7)kM#Ho_RWmiBp
RRRRnz4I:RRRRHV58IN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#Rp5BiW,Rq)772CRLo
HMRRRRRRRRRRRRH5VRBRpi=4R''MRN8pRBiP'CC2M0RC0EMR
RRRRRRRRRRRRRRNRI8C_so=R<R7Wq7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#S;
CRM8oCCMsCN0Rnz4IR;
RzRR4R(I:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);S8CMRMoCC0sNC4Rz(
I;
RRRRR-- sG0NFRDoRHOVRFs7DkNRsbF0NRO#SC
-7-RFFRM0CRMC08RERH#VRFsM8FsIEsO	NRO#-C
-sSzC:oRRFbsO#C#5iBp2CRLo
HM-R-SRRHV5iBp'  ehNaRMB8Rp=iRR''42ER0C-M
-RSRRh7Q_b0lRR<=7;Qh
S--R)RRq)77_b0lRR<=)7q7)-;
-RSRR7Wq70)_l<bR=qRW7;7)
S--RWRR l_0b=R<R;W 
S--RMRC8VRH;-
-S8CMRFbsO#C#;S

-Q-RVCR)Nq8R8C8s#=#RRHWs0qCR8C8s#R#,LN$b#7#RQ0hRFkRF00bkRRHVWH R#MRCNCLD8z
SlRkG:sRbF#OC#k5F0C_soS2
RCRLo
HM-R-SRHRRVWR5q)77_b0lR)=Rq)77_b0lR8NMR_W 0Rlb=4R''02RE
CM-S-SRkRF0C_so<4R=QR7hl_0b-;
-CSSD
#CSRSRF_k0s4CoRR<=F_k0s5CoI0H8ER-48MFI0jFR2-;
-CSSMH8RVS;
CRM8bOsFC;##
RSRRRR
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4__141S4
zR4U:VRHRE5OFCHO_8IH0=ERRR42oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RSRREzO	H:RVNR58I8sHE80R4>Rco2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24cRR<=)7q7)85N8HsI8-0E4FR8IFM0R24c;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SR8CMRMoCC0sNCORzE
	;RRRRSgz4RV:RFHsRRRHM5b8C0ME_kOl_C#DDR4-R2FR8IFM0RojRCsMCN
0CSR--Q5VRNs88I0H8ERR>4Rc2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRSRRzR.j:VRHR85N8HsI8R0E>cR42CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
SFSSkC0_M25HRR<='R4'IMECR_5sNs88_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=WI RERCM58IN_osC58N8s8IH04E-RI8FMR0F4Rc2=2RHR#CDCjR''R;
RRRRRSRRCRM8oCCMsCN0Rjz.;-
S-VRQR85N8HsI8R0E<4=RcM2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRSRRzRS.:4RRRHV58N8s8IH0<ER=cR42CRoMNCs0SC
SFSSkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;.4
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzR..:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq4v_ncdUXR47:NRDLRCDH"#RW
";RRRRRRRRRRRRRRRRLHCoMR
RRRRRRRRRRARS)_qv4Undc7X4R):Rq4vAn4_1_
14SRRRRRRRRRRRRsbF0NRlb7R5Qjq52>R=R_HMs5Co[R2,q)77q>R=RIDF_8IN84s5dFR8IFM0R,j2RA7QRR=>",j"R7q7)=AR>FRDIN_s858s48dRF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SRSSR7RRm=qR>bRFCRM,75mAj=2R>kRF0k_L#H45,2[2;R

RRRRRRRRRRRRRFRRks0_C[o52=R<R0Fk_#Lk4,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz.R;
RRRRS8CMRMoCC0sNC4RzgR;
RCRRMo8RCsMCNR0Cz;4URRRR
RRRR
RRRRRR-t-RCsMCNR0C0REC)RqvODCD#MRN8CR#D0CORoDFHVORF)sRq4vAn._1_
1.Sdz.RH:RVOR5EOFHCH_I8R0E=2R.RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
SREzO	RR:H5VRNs88I0H8ERR>4Rd2oCCMsCN0
RRRRRRRRDkO	RR:bOsFC5##B2pi
RRRRRRRRCRLo
HMRRRRRRRRRVRHRp5BiP'CCRM0NRM8BRpi=4R''02RE
CMRRRRRRRRRRRRs8_N8ss_CNo58I8sHE80-84RF0IMFdR42=R<R7)q7N)58I8sHE80-84RF0IMFdR42R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#RDkO	S;
RMRC8CRoMNCs0zCRO;E	
RRRR.SzcRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24dRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRS6z.RH:RVNR58I8sHE80R4>Rdo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24dRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNC.Rz6S;
-Q-RVNR58I8sHE80RR<=4Rd2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzR.n:VRHR85N8HsI8R0E<4=Rdo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNC.RznS;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRR.Sz(RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gU4.7X.RD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gU4.7X.R):Rq4vAn._1_
1.SRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[.*+84RF0IMF*R.[R2,q)77q>R=RIDF_8IN84s5.FR8IFM0R,j2RA7QRR=>""jj,7Rq7R)A=D>RFsI_Ns885R4.8MFI0jFR2S,
SRSRRhR q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SRSSR7RRm=qR>bRFCRM,75mA4=2R>kRF0k_L#H.5,[.*+,42RA7m5Rj2=F>RkL0_k5#.H.,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5.[<2R=kRF0k_L#H.5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C.o5*4[+2=R<R0Fk_#Lk.,5H.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNC.Rz(R;
RRRRS8CMRMoCC0sNC.RzcR;
RCRRMo8RCsMCNR0Cz;.dR
R
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_cc_1
.SzURR:H5VROHEFOIC_HE80Rc=R2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RORzER	:H5VRNs88I0H8ERR>4R.2oCCMsCN0RR
RRRRRRORkD:	RRFbsO#C#5iBp2R
RRRRRRLRRCMoH
RRRRRRRRHRRVBR5pCi'P0CMR8NMRiBpR'=R4R'20MEC
RRRRRRRRRRRRNs_8_8ss5CoNs88I0H8ER-48MFI04FR.<2R=qR)757)Ns88I0H8ER-48MFI04FR.
2;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#ORkD
	;SCRRMo8RCsMCNR0Cz	OE;R
RRzRS.:gRRsVFRHHRM8R5CEb0_lMk_DOCD-#RRR428MFI0jFRRMoCC0sNC-
S-VRQR85N8HsI8R0E>.R42CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdSzjRR:H5VRNs88I0H8ERR>4R.2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
RRRRRRRRRRRRRRRR0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RWRCIEMIR5Ns8_CNo58I8sHE80-84RF0IMF.R42RR=HC2RDR#C';j'
RRRRRRRRMSC8CRoMNCs0zCRd
j;SR--Q5VRNs88I0H8E=R<R24.RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
RRRRRS4zdRH:RVNR58I8sHE80RR<=4R.2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCdRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRdSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_gcjn7XcRD:RNDLCRRH#";W"
RRRRRRRRRRRRRRRRoLCHRM
RRRRRRRRRSRRAv)q_gcjn7XcR):Rq4vAnc_1_
1cSRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5[c*+8dRF0IMF*Rc[R2,q)77q>R=RIDF_8IN84s54FR8IFM0R,j2RA7QRR=>"jjjjR",q)77A>R=RIDF_8sN84s54FR8IFM0R,j2
SSSSq hRR=>',4'R)11q>R=R''j, RWq>R=R0Is_5CMHR2,BqpiRR=>B,piRA hRR=>',4'R)11A>R=R''j, RWA>R=R''j,pRBi=AR>pRBiS,
S7SSm=qR>bRFCRM,75mAd=2R>kRF0k_L#Hc5,*Rc[2+d,mR7A25.RR=>F_k0Lck#5cH,*.[+2
,RSSSS75mA4=2R>kRF0k_L#Hc5,[c*+,42RA7m5Rj2=F>RkL0_k5#cHc,R*2[2;R
RRRRRRRRRRRRRRkRF0C_so*5c[<2R=kRF0k_L#Hc5,[c*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cco5*4[+2=R<R0Fk_#Lkc,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Coc+*[.<2R=kRF0k_L#Hc5,[c*+R.2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[c*+Rd2<F=RkL0_k5#cH*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R

RRRRRSRRCRM8oCCMsCN0R.zd;R
RRSRRCRM8oCCMsCN0Rgz.;R
RRMRC8CRoMNCs0zCR.
U;
RSRR-R-RMtCC0sNCER0CqR)vCRODRD#NRM8#CCDOD0RFOoHRsVFRv)qA_4n11g_gz
Sd:dRRRHV5FOEH_OCI0H8ERR=go2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SzRRORE	:VRHR85N8HsI8R0E>4R42CRoMNCs0RC
RRRRRkRRORD	:sRbF#OC#p5BiR2
RRRRRRRRLHCoMR
RRRRRRRRRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMR
RRRRRRRRRR_RsNs88_osC58N8s8IH04E-RI8FMR0F4R42<)=Rq)7758N8s8IH04E-RI8FMR0F4;42
RRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#k#RO;D	
RSRCRM8oCCMsCN0REzO	R;
RSRRzRdc:FRVsRRHH5MR80CbEk_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0SC
-Q-RVNR58I8sHE80R4>R4M2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRRzRSd:6RRRHV58N8s8IH0>ERR244RMoCC0sNC-
S-HRVGFRVsNROD4DRd(UU,CR#D0CORRFV0#sH0CN0R0MFRHLCMsoRC#oH0CCs8R
RRRRRRRRRRRRRRkRF0M_C5RH2<'=R4I'RERCM5Ns_8_8ss5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R ERIC5MRI_N8s5CoNs88I0H8ER-48MFI04FR4=2RRRH2CCD#R''j;R
RRRRRRCRSMo8RCsMCNR0Cz;d6
-S-RRQV58N8s8IH0<ER=4R42FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
SRRRRdSznRR:H5VRNs88I0H8E=R<R244RMoCC0sNCR
SRRRRRRRRRFRRkC0_M25HRR<=';4'
RRRRRRRRRRRRRRRR0Is_5CMH<2R= RW;R
RRRRRRCRSMo8RCsMCNR0Cz;dn
-S-RMtCC0sNCER0CqR)vCRODRD#NRM80-sH#00NCR#
RRRRRSRRzRd(:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq.v_jXcUU:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
RRRRRRRRRRRR)SAq.v_jXcUU:7RRv)qA_4n11g_gR
RRRRRRRRRRRRRRRRRb0FsRblNRQ57q>R=R_HMs5Cog+*[(FR8IFM0R[g*2q,R7q7)RR=>D_FII8N8sj54RI8FMR0FjR2,7RQA=">Rjjjjjjjj"q,R7A7)RR=>D_FIs8N8sj54RI8FMR0Fj
2,SSSS Rhq='>R4R',1q1)RR=>',j'RqW RR=>I_s0CHM52B,RpRiq=B>RpRi, RhA='>R4R',1A1)RR=>',j'RAW RR=>',j'RiBpA>R=RiBp,SR
S7SSm=qR>bRFCRM,75mA(=2R>kRF0k_L#HU5,[U*+,(2RA7m5Rn2=F>RkL0_k5#UH*,U[2+n,SR
S7SSm6A52>R=R0Fk_#LkU,5HU+*[6R2,75mAc=2R>kRF0k_L#HU5,[U*+,c2RA7m5Rd2=F>RkL0_k5#UH*,U[2+d,SR
S7SSm.A52>R=R0Fk_#LkU,5HU+*[.R2,75mA4=2R>kRF0k_L#HU5,[U*+,42RA7m5Rj2=F>RkL0_k5#UH*,U[R2,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRu7Qq25jRR=>HsM_Cgo5*U[+27,RQRuA=">RjR",7qmuRR=>FMbC,mR7ujA52>R=RsbNH_0$LUk#5[H,2
2;RRRRRRRRRRRRRRRRF_k0s5Cog2*[RR<=F_k0LUk#5UH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R42<F=RkL0_k5#UH*,U[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+.RR<=F_k0LUk#5UH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*d[+2=R<R0Fk_#LkU,5HU+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[c<2R=kRF0k_L#HU5,[U*+Rc2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRRRRRR0Fk_osC5[g*+R62<F=RkL0_k5#UH*,U[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_so*5g[2+nRR<=F_k0LUk#5UH,*n[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_Cgo5*([+2=R<R0Fk_#LkU,5HU+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Cog+*[U<2R=NRbs$H0_#LkU,5H[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRS8CMRMoCC0sNCdRz(R;
RRRRS8CMRMoCC0sNCdRzcR;
RCRRMo8RCsMCNR0Cz;dd
R
SR-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOFRVsqR)vnA4_U14_U14
dSzURR:H5VROHEFOIC_HE80R4=RUo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8SRRRz	OERH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CRRRRRRRRk	ODRb:RsCFO#B#5p
i2RRRRRRRRRoLCHRM
RRRRRRRRRRHV5iBp'CCPMN0RMB8Rp=iRR''42ER0CRM
RRRRRRRRRsRR_8N8sC_so85N8HsI8-0E4FR8IFM0R24jRR<=)7q7)85N8HsI8-0E4FR8IFM0R24j;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFCR##k	OD;R
SRMRC8CRoMNCs0zCRO;E	
RRRRdSzgRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERR24jRCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRSjzcRH:RVNR58I8sHE80R4>Rjo2RCsMCN
0CSR--VRHGVRFsODNDRU4dUR(,#CCDOF0RVsR0HN#00MCRFL0RCoHMRosCHC#0s
C8RRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5_8N8sC_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0R24jRH=R2DRC#'CRj
';RRRRRRRRS8CMRMoCC0sNCcRzjS;
-Q-RVNR58I8sHE80RR<=4Rj2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRSRSRRzRc4:VRHR85N8HsI8R0E<4=Rjo2RCsMCN
0CSRRRRRRRRRRRR0Fk_5CMH<2R=4R''R;
RRRRRRRRRRRRRIRRsC0_M25HRR<=W
 ;RRRRRRRRS8CMRMoCC0sNCcRz4S;
-t-RCsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcSz.RR:VRFs[MRHRH5I8_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVAv)q_.4jcnX47RR:DCNLD#RHR""W;R
RRRRRRRRRRRRRRCRLo
HMRRRRRRRRRRRRSqA)vj_4.4cXn:7RRv)qA_4n1_4U1
4URRRRRRRRRRRRRRRRRFRbsl0RN5bR7RQq=H>RMC_soU54*4[+6FR8IFM0R*4U[R2,q)77q>R=RIDF_8IN8gs5RI8FMR0FjR2,7RQA=">Rjjjjjjjjjjjjjjjj"q,R7A7)RR=>D_FIs8N8sR5g8MFI0jFR2S,
S SSh=qR>4R''1,R1R)q='>RjR',WR q=I>RsC0_M25H,pRBi=qR>pRBi ,Rh=AR>4R''1,R1R)A='>RjR',WR A='>RjR',BApiRR=>B,piRS
SSmS7q>R=RCFbM7,Rm4A56=2R>kRF0k_L#54nHn,4*4[+6R2,75mA4Rc2=F>RkL0_kn#454H,n+*[4,c2RS
SSmS7Ad542>R=R0Fk_#Lk4Hn5,*4n[d+427,Rm4A5.=2R>kRF0k_L#54nHn,4*4[+.R2,75mA4R42=F>RkL0_kn#454H,n+*[4,42RS
SSmS7Aj542>R=R0Fk_#Lk4Hn5,*4n[j+427,RmgA52>R=R0Fk_#Lk4Hn5,*4n[2+g,mR7A25URR=>F_k0L4k#n,5H4[n*+,U2RS
SSmS7A25(RR=>F_k0L4k#n,5H4[n*+,(2RA7m5Rn2=F>RkL0_kn#454H,n+*[nR2,75mA6=2R>kRF0k_L#54nHn,4*6[+2
,RSSSS75mAc=2R>kRF0k_L#54nHn,4*c[+27,RmdA52>R=R0Fk_#Lk4Hn5,*4n[2+d,mR7A25.RR=>F_k0L4k#n,5H4[n*+,.2RS
SSmS7A254RR=>F_k0L4k#n,5H4[n*+,42RA7m5Rj2=F>RkL0_kn#454H,n2*[,RR
RRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_soU54*4[+(FR8IFM0R*4U[n+427,RQRuA=">Rj,j"Ru7mq>R=RCFbMR,
RRRRRRRRRRRRRRRRRRRRRRRRR7RRm5uA4=2R>NRbs$H0_#Lk4Hn5,[.*+,42Ru7mA25jRR=>bHNs0L$_kn#45.H,*2[2;R
RRRRRRRRRRRRRRkRF0C_soU54*R[2<F=RkL0_kn#454H,n2*[RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+2=R<R0Fk_#Lk4Hn5,*4n[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*.[+2=R<R0Fk_#Lk4Hn5,*4n[2+.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*d[+2=R<R0Fk_#Lk4Hn5,*4n[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*c[+2=R<R0Fk_#Lk4Hn5,*4n[2+cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*6[+2=R<R0Fk_#Lk4Hn5,*4n[2+6RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*n[+2=R<R0Fk_#Lk4Hn5,*4n[2+nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*([+2=R<R0Fk_#Lk4Hn5,*4n[2+(RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*U[+2=R<R0Fk_#Lk4Hn5,*4n[2+URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*g[+2=R<R0Fk_#Lk4Hn5,*4n[2+gRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+j<2R=kRF0k_L#54nHn,4*4[+jI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+244RR<=F_k0L4k#n,5H4[n*+244RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+.<2R=kRF0k_L#54nHn,4*4[+.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+24dRR<=F_k0L4k#n,5H4[n*+24dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+c<2R=kRF0k_L#54nHn,4*4[+cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';RRRRRRRRRRRRRRRRF_k0s5Co4[U*+246RR<=F_k0L4k#n,5H4[n*+246RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRRRRRRRRRkRF0C_soU54*4[+n<2R=NRbs$H0_#Lk4Hn5,[.*2ERIC5MRF_k0CHM52RR='24'R#CDCZR''R;
RRRRRRRRRRRRRFRRks0_C4o5U+*[4R(2<b=RN0sH$k_L#54nH*,.[2+4RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;R
RRRRRRCRSMo8RCsMCNR0Cz;c.
RRRRCRSMo8RCsMCNR0Cz;dg
RRRR8CMRMoCC0sNCdRzU
;
SRRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDoRHOVRFs)Aqv41n_d1n_dSn
zNdURH:RVOR5EOFHCH_I8R0E=nRd2CRoMNCs0SC
-V-RHVGRFOsRNRDD4UdU(#,RCODC0VRFRH0s#00NCFRM0CRLHRMosHCo#s0CCS8
RzRRORE	:VRHR85N8HsI8R0E>2RgRMoCC0sNCR
SRkRRORD	:sRbF#OC#p5BiS2
SCRLo
HMSRSRH5VRB'piCMPC0MRN8pRBiRR='24'RC0EMS
SRRRRs8_N8ss_CNo58I8sHE80-84RF0IMF2RgRR<=)7q7)85N8HsI8-0E4FR8IFM0R;g2
RSSR8CMR;HV
CSSMb8RsCFO#k#RO;D	
RSRR8CMRMoCC0sNCORzE
	;SRRRRgzdNRR:VRFsHMRHRC58b_0EM_klODCD#RR-482RF0IMFRRjoCCMsCN0
-S-RRQV58N8s8IH0>ERRRg2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHSO
ScSzj:NRRRHV58N8s8IH0>ERRRg2oCCMsCN0
-S-RGVHRsVFRDONDdR4U,U(RD#CCRO0F0VRs0H#NR0CMRF0LMCHoCRso0H#C8sC
SSSS0Fk_5CMH<2R=4R''ERIC5MRs8_N8ss_CNo58I8sHE80-84RF0IMF2RgRH=R2DRC#'CRj
';SSSSI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRg2=2RHR#CDCjR''S;
SMSC8CRoMNCs0zCRc;jN
-S-RRQV58N8s8IH0<ER=2RgRRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88S
SS4zcNRR:H5VRNs88I0H8E=R<RRg2oCCMsCN0
SSSS0Fk_5CMH<2R=4R''S;
SISSsC0_M25HRR<=W
 ;SCSSMo8RCsMCNR0CzNc4;-
S-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#SzSScR.N:FRVsRR[H5MRI0H8Ek_MlC_ODRD#-2R4RI8FMR0FjCRoMNCs0RC
RRRRRRRRRRRRRNRR0H0sLCk0Rs\3NFl_VCV#0F\RV)RAq6v_4d.X.:7RRLDNCHDR#WR""R;
RRRRRRRRRRRRRLRRCMoH
SSSSqA)v4_6..Xd7RR:)Aqv41n_d1n_dRn
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsbF0NRlb7R5Q=qR>MRH_osC5*dn[4+dRI8FMR0Fd[n*2q,R7q7)RR=>D_FII8N8sR5U8MFI0jFR27,RQ=AR>jR"jjjjjjjjjjjjjjjjjjjjjjjjjjjjj"jj,7Rq7R)A=D>RFsI_Ns8858URF0IMF2Rj,S
SShS q>R=R''4,1R1)=qR>jR''W,R =qR>sRI0M_C5,H2RiBpq>R=RiBp,hR A>R=R''4,1R1)=AR>jR''W,R =AR>jR''B,RpRiA=B>Rp
i,SSSS7Rmq=F>Rb,CMRA7m52d4RR=>F_k0Ldk#.,5Hd[.*+2d4,mR7Aj5d2>R=R0Fk_#LkdH.5,*d.[j+d2S,
S7SSm.A5g=2R>kRF0k_L#5d.H.,d*.[+gR2,75mA.RU2=F>RkL0_k.#d5dH,.+*[.,U2RA7m52.(RR=>F_k0Ldk#.,5Hd[.*+2.(,S
SSmS7An5.2>R=R0Fk_#LkdH.5,*d.[n+.27,Rm.A56=2R>kRF0k_L#5d.H.,d*.[+6R2,75mA.Rc2=F>RkL0_k.#d5dH,.+*[.,c2
SSSSA7m52.dRR=>F_k0Ldk#.,5Hd[.*+2.d,mR7A.5.2>R=R0Fk_#LkdH.5,*d.[.+.27,Rm.A54=2R>kRF0k_L#5d.H.,d*.[+4
2,SSSS75mA.Rj2=F>RkL0_k.#d5dH,.+*[.,j2RA7m524gRR=>F_k0Ldk#.,5Hd[.*+24g,mR7AU542>R=R0Fk_#LkdH.5,*d.[U+42S,
S7SSm4A5(=2R>kRF0k_L#5d.H.,d*4[+(R2,75mA4Rn2=F>RkL0_k.#d5dH,.+*[4,n2RA7m5246RR=>F_k0Ldk#.,5Hd[.*+246,S
SSmS7Ac542>R=R0Fk_#LkdH.5,*d.[c+427,Rm4A5d=2R>kRF0k_L#5d.H.,d*4[+dR2,75mA4R.2=F>RkL0_k.#d5dH,.+*[4,.2
SSSSA7m5244RR=>F_k0Ldk#.,5Hd[.*+244,mR7Aj542>R=R0Fk_#LkdH.5,*d.[j+427,RmgA52>R=R0Fk_#LkdH.5,*d.[2+g,S
SSmS7A25URR=>F_k0Ldk#.,5Hd[.*+,U2RA7m5R(2=F>RkL0_k.#d5dH,.+*[(R2,75mAn=2R>kRF0k_L#5d.H.,d*n[+2S,
S7SSm6A52>R=R0Fk_#LkdH.5,*d.[2+6,mR7A25cRR=>F_k0Ldk#.,5Hd[.*+,c2RA7m5Rd2=F>RkL0_k.#d5dH,.+*[d
2,SSSS75mA.=2R>kRF0k_L#5d.H.,d*.[+27,Rm4A52>R=R0Fk_#LkdH.5,*d.[2+4,mR7A25jRR=>F_k0Ldk#.,5Hd[.*2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR7RRQRuq=H>RMC_son5d*d[+6FR8IFM0R*dn[.+d27,RQRuA=">Rjjjj"7,RmRuq=F>Rb,CM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA25dRR=>bHNs0L$_k.#d5cH,*d[+27,Rm5uA.=2R>NRbs$H0_#LkdH.5,[c*+,.2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRu7mA254RR=>bHNs0L$_k.#d5cH,*4[+27,Rm5uAj=2R>NRbs$H0_#LkdH.5,[c*2
2;SSSSF_k0s5Cod[n*2=R<R0Fk_#LkdH.5,*d.[I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+R42<F=RkL0_k.#d5dH,.+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+R.2<F=RkL0_k.#d5dH,.+*[.I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+Rd2<F=RkL0_k.#d5dH,.+*[dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+Rc2<F=RkL0_k.#d5dH,.+*[cI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+R62<F=RkL0_k.#d5dH,.+*[6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+Rn2<F=RkL0_k.#d5dH,.+*[nI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+R(2<F=RkL0_k.#d5dH,.+*[(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+RU2<F=RkL0_k.#d5dH,.+*[UI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+Rg2<F=RkL0_k.#d5dH,.+*[gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24jRR<=F_k0Ldk#.,5Hd[.*+24jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+4<2R=kRF0k_L#5d.H.,d*4[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24.RR<=F_k0Ldk#.,5Hd[.*+24.RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+d<2R=kRF0k_L#5d.H.,d*4[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24cRR<=F_k0Ldk#.,5Hd[.*+24cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+6<2R=kRF0k_L#5d.H.,d*4[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24nRR<=F_k0Ldk#.,5Hd[.*+24nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+(<2R=kRF0k_L#5d.H.,d*4[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+24URR<=F_k0Ldk#.,5Hd[.*+24URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*4[+g<2R=kRF0k_L#5d.H.,d*4[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.jRR<=F_k0Ldk#.,5Hd[.*+2.jRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+4<2R=kRF0k_L#5d.H.,d*.[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2..RR<=F_k0Ldk#.,5Hd[.*+2..RCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+d<2R=kRF0k_L#5d.H.,d*.[+dI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.cRR<=F_k0Ldk#.,5Hd[.*+2.cRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+6<2R=kRF0k_L#5d.H.,d*.[+6I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.nRR<=F_k0Ldk#.,5Hd[.*+2.nRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+(<2R=kRF0k_L#5d.H.,d*.[+(I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2.URR<=F_k0Ldk#.,5Hd[.*+2.URCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*.[+g<2R=kRF0k_L#5d.H.,d*.[+gI2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2djRR<=F_k0Ldk#.,5Hd[.*+2djRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SSkSF0C_son5d*d[+4<2R=kRF0k_L#5d.H.,d*d[+4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2d.RR<=bHNs0L$_k.#d5cH,*R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
SSSS0Fk_osC5*dn[d+d2=R<RsbNH_0$Ldk#.,5Hc+*[4I2RERCM50Fk_5CMH=2RR''42DRC#'CRZ
';SSSSF_k0s5Cod[n*+2dcRR<=bHNs0L$_k.#d5cH,*.[+2ERIC5MRF_k0CHM52RR='24'R#CDCZR''S;
SFSSks0_Cdo5n+*[dR62<b=RN0sH$k_L#5d.H*,c[2+dRCIEMFR5kC0_M25HR'=R4R'2CCD#R''Z;S
SS8CMRMoCC0sNCcRz.
N;SMSC8CRoMNCs0zCRd;gN
MSC8CRoMNCs0zCRd;UN
CRRMo8RCsMCNR0Cz;cd
R
RzRcc:VRHRF5M0NRs8_8ss2CoRMoCC0sNC-R-RMoCC0sNCCR#D0CORlsN
RRRRR--QNVR8I8sHE80R6<RR#N#HRoM'Rj'0kFRMCk#8HRL0R#
RzRRj:RRRRHV58N8s8IH0=ERRR42oCCMsCN0
RRRRRRRRIDF_8sN8#s_RR<="jjjjRj"&NRs8C_so5_#j
2;RRRRRRRRD_FII8N8sR_#<"=Rjjjjj&"RR8IN_osC_j#52R;
RCRRMo8RCsMCNR0Cz
j;RRRRzR4R:VRHR85N8HsI8R0E=2R.RMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"jjRj"&NRs8C_so5_#4FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<="jjjj&"RR8IN_osC_4#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;z4
RRRRRz.RH:RVNR58I8sHE80Rd=R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=jR"jRj"&NRs8C_so5_#.FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<="jjj"RR&I_N8s_Co#R5.8MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RcRMoCC0sNCR
RRRRRRFRDIN_s8_8s#=R<Rj"j"RR&s_N8s_Co#R5d8MFI0jFR2R;
RRRRRDRRFII_Ns88_<#R=jR"j&"RR8IN_osC_d#5RI8FMR0Fj
2;RRRRCRM8oCCMsCN0R;zd
cSzSH:RVNR58I8sHE80R6=R2CRoMNCs0SC
SIDF_8sN8#s_RR<='Rj'&NRs8C_so5_#cFR8IFM0R;j2
DSSFII_Ns88_<#R=jR''RR&I_N8s_Co#R5c8MFI0jFR2S;
CRM8oCCMsCN0R;zc
RRRRRz6RH:RVNR58I8sHE80R6>R2CRoMNCs0RC
RRRRRDRRFsI_Ns88_<#R=NRs8C_so5_#6FR8IFM0R;j2
RRRRRRRRIDF_8IN8#s_RR<=I_N8s_Co#R568MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
6;
RRRRR--Q5VR8_HMs2CoRosCHC#0sQR7h#RkHRMoB
piRRRRzRnR:VRHRH58MC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,QR7hL2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRHRRMC_soR_#<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNCnRz;R
RR(RzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osC_<#R=QR7hR;
RCRRMo8RCsMCNR0Cz
(;
RRRRR--Q5VR80Fk_osC2CRso0H#C7sRmRzakM#HoBRmpRi
RzRRU:RRRRHV5k8F0C_soo2RCsMCN
0CRRRRRRRRbOsFCR##5pmBiF,Rks0_C#o_2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s_Co#R;
RRRRRRRRRCRRMH8RVR;
RRRRRCRRMb8RsCFO#
#;RRRRCRM8oCCMsCN0R;zU
RRRRRzgRH:RVMR5F80RF_k0s2CoRMoCC0sNCR
RRRRRRRRRRmR7z<aR=kRF0C_so;_#
RRRR8CMRMoCC0sNCgRz;R

R-RR-VRQR85N8ss_CRo2sHCo#s0CR7q7)#RkHRMoB
piRRRRzR4jRH:RVsR5Ns88_osC2CRoMNCs0RC
RRRRRbRRsCFO#5#RB,piR7)q7R)2LHCoMR
RRRRRRRRRRVRHRp5BiRR='R4'NRM8B'piCMPC002RE
CMRRRRRRRRRRRRRRRRs_N8s_Co#=R<R7)q7N)58I8sHE80-84RF0IMF2Rj;R
RRRRRRRRRRMRC8VRH;R
RRRRRRMRC8sRbF#OC#R;
RCRRMo8RCsMCNR0Cz;4j
RRRR4z4RH:RVMR5Fs0RNs88_osC2CRoMNCs0RC
RRRRRRRRRsRRNs8_C#o_RR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;44
R
RR-R-RRQV58N8sC_sos2RC#oH0RCsq)77RHk#MBoRpRi
RzRR4R.R:VRHRN5I8_8ss2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,W7q7)L2RCMoH
RRRRRRRRRRRRRHV5iBpR'=R4N'RMB8RpCi'P0CM2ER0CRM
RRRRRRRRRRRRRIRRNs8_C#o_RR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
.;RRRRzR4d:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_soR_#<W=Rq)77;R
RRMRC8CRoMNCs0zCR4
d;RRRRRRRR
RRRRR--tCCMsCN0RC0ERv)qRDOCDN#RM#8RCODC0FRDo
HORRRRzR4c:FRVsRRHH5MRM_klODCD_Rnc-2R4RI8FMR0FjCRoMNCs0RC
R-RR-VRQR85N8HsI8R0E>2R6RCMC8FR0RCOsNR0CI0sHCMRCNCLDR8NMR0FkbRk0CLMND#CRCODC0FRDo
HORRRRRRRRzR46:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_H#52=R<R''4RCIEMsR5Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRRH2CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_H#52=R<RRW IMECRN5I8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=HC2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC4Rz6R;
R-RR-VRQR85N8HsI8R0E<6=R2FRMRHIs0CCRMDNLCsRFR0FkbRk0CLMND#CRCODC0FRDoRHOM8CCCR8
RRRRRzRR4:nRRRHV58N8s8IH0<ER=2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_H#52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C_H#52=R<R;W 
RRRRRRRR8CMRMoCC0sNC4RznR;
R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRH0s-N#00
C#RRRRRRRRzR4(:FRVsRR[H5MRI0H8ERR-482RF0IMFRRjoCCMsCN0
RRRRRRRRRRRR0N0skHL0\CR3lsN_VFV#\C0RRFVzv)qn:cRRLDNCHDR#1R"7Ra"&MRH0CCosl'HN5oCI0H8E&2RR""7RH&RMo0CCHs'lCNo5nH*c&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50E54H+2c*n,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qn:cRRqX)vXnc4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,q=6R>FRDIN_I8_8s#256,SR
SSSSS7RRuj)qRR=>D_FIs8N8s5_#jR2,7qu)4>R=RIDF_8sN8#s_5,42R)7uq=.R>FRDIN_s8_8s#25.,S
SSSSSRuR7)Rqd=D>RFsI_Ns88_d#527,Ruc)qRR=>D_FIs8N8s5_#cR2,7qu)6>R=RIDF_8sN8#s_5,62RS
SSSSSR RWRR=>I_s0C#M_5,H2RpWBi>R=RiBp,uR7m>R=R0Fk_#Lk_#nc5[H,2
2;RRRRRRRRRRRRRRRRF_k0s_Co#25[RR<=F_k0L_k#n5c#H2,[RCIEMFR5kC0_M5_#H=2RR''42DRC#'CRZ
';RRRRRRRRCRM8oCCMsCN0R(z4;R
RRCRRMo8RCsMCNR0Cz;4cRRRRRRRRRRRR
RRRR
RRRRRR-t-RCsMCNR0CN.RdRsIF8CR8C)bRqOvRCRDDHNVRbFbsbNsH0RCRRRRRRRRRRRRRRR
RR4RzURR:H5VRM_klODCD_Rd.=2R4RMoCC0sNCR
RR-R-RRQV58N8s8IH0>ERRR(2M8CCRR0FONsC0ICRsCH0RNCMLRDCNRM8Fbk0kC0RMDNLCCR#D0CORoDFHRO
RRRRRzRR4RgN:VRHR85N8HsI8R0E>2RnRMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_Rd.<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''j2C2RDR#C';j'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RWRCIEM5R5I_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58RI_N8s_Co#256R'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN4g;R
RRRRRR4Rzg:LRRRHV58N8s8IH0=ERRNnRMM8RkOl_C_DDn=cRRRj2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CMd<.R=4R''ERIC5MR58sN_osC_6#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CdM_.=R<RRW IMECRI55Ns8_C#o_5R62=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR4;gLRRRR-Q-RVNR58I8sHE80RR<=6M2RFsRIHR0CCLMNDFCRskRF00bkRNCMLRDC#CCDOD0RFOoHRCMC8
C8RRRRRRRRzR.j:VRHR85N8HsI8R0E<6=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_M._dRR<=';4'
RRRRRRRRRRRRRRRR0Is__CMd<.R= RW;R
RRRRRRMRC8CRoMNCs0zCR.
j;RRRR-t-RCsMCNR0C0REC)RqvODCDR8NMRH0s-N#00RC
RRRRRzRR.:4RRsVFRH[RMIR5HE80R4-R2FR8IFM0RojRCsMCN
0CRRRRRRRRRRRRNs00H0LkC3R\s_NlF#VVCR0\FzVR)dqv.RR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCM_klODCD_*ncnRc2&WR""RR&HCM0o'CsHolNC25[R"&R &"RR0HMCsoC'NHlooC5CC0_M88_CEb05lMk_DOCDc_n*Rnc+.Rd,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)qd:.RRqX)vXd.4
7RRRRRRRRRRRRRRRRRb0FsRblNRR57=H>RMC_so5_#[R2,q=jR>FRDIN_I8_8s#25j,4RqRR=>D_FII8N8s5_#4R2,q=.R>FRDIN_I8_8s#25.,R
RRRRRRRRRRRRRRRRRRRRRRRRRq=dR>FRDIN_I8_8s#25d,cRqRR=>D_FII8N8s5_#cR2,
SSSSRSSR)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2R)7uq=cR>FRDIN_s8_8s#25c,SR
SSSSSWRR >R=R0Is__CMdR.,WiBpRR=>B,piRm7uRR=>F_k0L_k#d5.#M_klODCD_,d.[;22
RRRRRRRRRRRRRRRR0Fk_osC_[#52=R<R0Fk_#Lk_#d.5lMk_DOCD._d,R[2IMECRk5F0M_C_Rd.=4R''C2RDR#C';Z'
RRRRRRRRMRC8CRoMNCs0zCR.
4;RRRRR8CMRMoCC0sNC4RzUR;RRRRRRRRR
R
RR-R-RMtCC0sNCRRN4InRFRs88bCCRv)qRDOCDVRHRbNbssFbHCN0RRRRRRRRRRRRR
RRRRRRzR..:VRHRk5MlC_OD4D_nRR=4o2RCsMCN
0CRRRR-Q-RVNR58I8sHE80R6>R2CRMC08RFsROCCN0RHIs0CCRMDNLCMRN8kRF00bkRNCMLRDC#CCDOD0RFOoH
RRRRRRRRdz.NRR:H5VRNs88I0H8ERR>nMRN8kRMlC_ODdD_.RR=4o2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0C4M_n=R<R''4RCIEM5R5s_N8s_Co#85N8HsI8-0E4FR8IFM0RRn2=kRMlC_ODnD_cN2RM58Rs_N8s_Co#256R'=R4R'2NRM858sN_osC_c#52RR='2j'2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0C4M_n=R<RRW IMECRI55Ns8_C#o_58N8s8IH04E-RI8FMR0Fn=2RRlMk_DOCDc_n2MRN8IR5Ns8_C#o_5R62=4R''N2RM58RI_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRCRRMo8RCsMCNR0CzN.d;R
RRRRRR.Rzd:LRRRHV58N8s8IH0>ERRNnRMM8RkOl_C_DDd/.R=2R4RMoCC0sNCR
RRRRRRRRRRRRRRkRF0M_C_R4n<'=R4I'RERCM5N5s8C_so5_#Ns88I0H8ER-48MFI0nFR2RR=M_klODCD_2ncR8NMRN5s8C_so5_#6=2RR''j2MRN8sR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRRRRRRRRRsRI0M_C_R4n<W=R ERIC5MR58IN_osC_N#58I8sHE80-84RF0IMF2RnRM=RkOl_C_DDnRc2NRM858IN_osC_6#52RR='2j'R8NMRN5I8C_so5_#c=2RR''j2C2RDR#C';j'
RRRRRRRR8CMRMoCC0sNC.Rzd
L;RRRRRRRRzO.dRH:RVNR58I8sHE80Rn=RR8NMRlMk_DOCD._dR4=R2CRoMNCs0RC
RRRRRRRRRRRRRFRRkC0_Mn_4RR<='R4'IMECRs55Ns8_C#o_5R62=4R''N2RM58Rs_N8s_Co#25cR'=Rj2'2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#6=2RR''42MRN8IR5Ns8_C#o_5Rc2=jR''R22CCD#R''j;R
RRRRRRMRC8CRoMNCs0zCR.;dO
RRRRRRRRdz.8RR:H5VRNs88I0H8ERR=6MRN8kRMlC_ODdD_.=R/RR42oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''ERIC5MR58sN_osC_N#58I8sHE80-84RF0IMF2RcRM=RkOl_C_DDd2.2R#CDCjR''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=WI RERCM5N5I8C_so5_#Ns88I0H8ER-48MFI0cFR2RR=M_klODCD_2d.2DRC#'CRj
';RRRRRRRRCRM8oCCMsCN0Rdz.8R;RR-R-RRQV58N8s8IH0<ER=2R6RRMFI0sHCMRCNCLDRRFsFbk0kC0RMDNLCCR#D0CORoDFHMORCCC88R
RRRRRR.RzcRR:H5VRNs88I0H8E=R<RRc2oCCMsCN0
RRRRRRRRRRRRRRRR0Fk__CM4<nR=4R''R;
RRRRRRRRRRRRRIRRsC0_Mn_4RR<=W
 ;RRRRRRRRCRM8oCCMsCN0Rcz.;R
RR-R-RMtCC0sNCER0CqR)vCRODNDRM08Rs#H-0CN0
RRRRRRRR6z.RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vR4n:NRDLRCDH"#R1"7aRH&RMo0CCHs'lCNo58IH0RE2&7R""RR&HCM0o'CsHolNCk5MlC_ODnD_cc*nRM+RkOl_C_DDdd.*.&2RR""WRH&RMo0CCHs'lCNo5R[2& R""RR&HCM0o'CsHolNCC5o0M_C8C_8b50EM_klODCD_*ncn+cRRlMk_DOCD._d*Rd.+nR4,CR8b20E2RR&"RX"&MRH0CCosl'HN5oC[2+4;R
RRRRRRRRRRCRLo
HMRRRRRRRRRRRRzv)q4:nRRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC_[#52q,Rj>R=RIDF_8IN8#s_5,j2RRq4=D>RFII_Ns88_4#52q,R.>R=RIDF_8IN8#s_5,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8#s_5,d2R)7uq=jR>FRDIN_s8_8s#25j,uR7)Rq4=D>RFsI_Ns88_4#527,Ru.)qRR=>D_FIs8N8s5_#.
2,SSSSSRSR7qu)d>R=RIDF_8sN8#s_5,d2RRW =I>RsC0_Mn_4,BRWp=iR>pRBi7,Ru=mR>kRF0k_L#n_4#k5MlC_OD4D_n2,[2R;
RRRRRRRRRRRRRFRRks0_C#o_5R[2<F=RkL0_k4#_nM#5kOl_C_DD4[n,2ERIC5MRF_k0C4M_nRR='24'R#CDCZR''R;
RRRRRCRRMo8RCsMCNR0Cz;.6
RRRR8CMRMoCC0sNC.Rz.R;RRRR
R8CMRMoCC0sNCcRzcC;
MN8RsHOE00COkRsCMsF_IE_OC;O	
-
-
R--p0N#RbHlDCClM00NHRFMH8#RCkVND-0
-s
NO0EHCkO0s#CRCODC0N_slVRFRv)q_W)_R
H#VOkM0MHFR0oC_8CM_b8C0#E5HRxC:MRH0CCosRR;80CbERR:HCM0o2CsR0sCkRsMHCM0oRCsHP#
NNsHLRDCl_HM#CHxRH:RMo0CC:sR=;Rj
oLCHRM
RMlH_x#HC=R:Rb8C0
E;RVRHRH5#x<CRRb8C0RE20MEC
RRRRMlH_x#HC=R:Rx#HCR;
R8CMR;HV
sRRCs0kMHRlMH_#x
C;CRM8o_C0C_M880CbEO;
F0M#NRM0M_klODCD#RR:HCM0oRCs:5=R5b8C0-ERR/424;n2RRRRRRRRRRRR-y-RRRFV)4qvn7X4RDOCDM#RCCC88$
0bFCRkL0_k0#_$RbCHN#Rs$sNRk5MlC_ODRD#8MFI0jFR,HRI8-0E4FR8IFM0RRj2F#VR0D8_FOoH;H
#oDMNR0Fk_#LkRF:RkL0_k0#_$;bCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-7R.RsNsNF$RVFR8k50RHkMb0FR0RH0s-N#002C#
o#HMRNDF_k0C:MRR8#0_oDFHPO_CFO0sk5MlC_ODRD#8MFI0jFR2R;RRRRRR-R-RNCML#DCRsVFRH0s-N#00
C##MHoNIDRsC0_MRR:#_08DHFoOC_POs0F5lMk_DOCD8#RF0IMF2Rj;RRRRRRRRR--I0sHCMRCNCLD#FRVsNRCOsERFFIRVqR)vCROD
D##MHoNHDRMC_soRR:#_08DHFoOC_POs0F58IH04E-RI8FMR0FjR2;RRRRRRRRRR--k8#CRR0FsHCo#s0CRh7QRH
#oDMNR0Fk_osCR#:R0D8_FOoH_OPC05FsI0H8ER-48MFI0jFR2R;RRRRRR-RR-#RkC08RFCRso0H#C7sRm
za#MHoNsDRNs8_C:oRR8#0_oDFHPO_CFO0s85N8HsI8-0E4FR8IFM0R;j2RRRRRR--k8#CRR0FsHCo#s0CR7)q7#)
HNoMDNRI8C_soRR:#_08DHFoOC_POs0F58N8s8IH04E-RI8FMR0FjR2;RRRR-k-R#RC80sFRC#oH0RCsW7q7)H
#oDMNRIDF_8sN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRs8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC2H
#oDMNRIDF_8IN8:sRR8#0_oDFHPO_CFO0sR5d8MFI0jFR2R;RRRRRRRRRR-RR-NRI8R8sL#H0RbHMk00RFqR)vCRODRD#5LcRHR0#skCJH8sC20
N0LsHkR0C\N3slV_FV0#C\RR:#H0sM
o;
oLCH
M
RRRR-Q-RV8RN8HsI8R0E<RRcNH##o'MRj0'RFMRkk8#CR0LH#R
RR4RzRRR:H5VRNs88I0H8ERR=4o2RCsMCN
0CRRRRRRRRD_FIs8N8s=R<Rj"jj&"RR8sN_osC5;j2
RRRRRRRRIDF_8IN8<sR=jR"jRj"&NRI8C_so25j;R
RRMRC8CRoMNCs0zCR4R;
RzRR.:RRRRHV58N8s8IH0=ERRR.2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=jR"j&"RR8sN_osC584RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<"=RjRj"&NRI8C_soR548MFI0jFR2R;
RCRRMo8RCsMCNR0Cz
.;RRRRzRdR:VRHR85N8HsI8R0E=2RdRMoCC0sNCR
RRRRRRFRDIN_s8R8s<'=Rj&'RR8sN_osC58.RF0IMF2Rj;R
RRRRRRFRDIN_I8R8s<'=Rj&'RR8IN_osC58.RF0IMF2Rj;R
RRMRC8CRoMNCs0zCRdR;
RzRRc:RRRRHV58N8s8IH0>ERRRd2oCCMsCN0
RRRRRRRRIDF_8sN8<sR=NRs8C_soR5d8MFI0jFR2R;
RRRRRDRRFII_Ns88RR<=I_N8s5CodFR8IFM0R;j2
RRRR8CMRMoCC0sNCcRz;R

R-RR-VRQRH58MC_sos2RC#oH0RCs7RQhkM#HopRBiR
RR6RzRRR:H5VR8_HMs2CoRMoCC0sNCR
RRRRRRsRbF#OC#BR5pRi,72QhRoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR_HMsRCo<7=RQ
h;RRRRRRRRRRRRCRM8H
V;RRRRRRRRCRM8bOsFC;##
RRRR8CMRMoCC0sNC6Rz;R
RRnRzRRR:H5VRMRF08_HMs2CoRMoCC0sNCR
RRRRRRRRRRMRH_osCRR<=7;Qh
RRRR8CMRMoCC0sNCnRz;R

R-RR-VRQRF58ks0_CRo2sHCo#s0CRz7ma#RkHRMomiBp
RRRRRz(RH:RV8R5F_k0s2CoRMoCC0sNCR
RRRRRRsRbF#OC#mR5B,piR0Fk_osC2CRLo
HMRRRRRRRRRRRRH5VRmiBpR'=R4N'RMm8RB'piCMPC002RE
CMRRRRRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR(R;
RzRRU:RRRRHV50MFRk8F0C_soo2RCsMCN
0CRRRRRRRRRRRR7amzRR<=F_k0s;Co
RRRR8CMRMoCC0sNCURz;R

R-RR-VRQRN5s8_8ss2CoRosCHC#0sqR)7R7)kM#HoBRmpRi
RzRRg:RRRRHV58sN8ss_CRo2oCCMsCN0
RRRRRRRRFbsO#C#RB5mpRi,)7q7)L2RCMoH
RRRRRRRRRRRRRHV5pmBiRR='R4'NRM8miBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8sN_osCRR<=)7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCRgR;
RzRR4:jRRRHV50MFR8sN8ss_CRo2oCCMsCN0
RRRRRRRRRRRR8sN_osCRR<=)7q7)R;
RCRRMo8RCsMCNR0Cz;4j
RRRRRRRRR
RR-R-RRQV58IN8ss_CRo2sHCo#s0CR7Wq7k)R#oHMRiBp
RRRR6z4RRR:H5VRI8N8sC_soo2RCsMCN
0CRRRRRRRRbOsFCR##5iBp,qRW727)RoLCHRM
RRRRRRRRRHRRVBR5p=iRR''4R8NMRiBp'CCPMR020MEC
RRRRRRRRRRRRRRRR8IN_osCRR<=W7q7)85N8HsI8-0E4FR8IFM0R;j2
RRRRRRRRRRRR8CMR;HV
RRRRRRRR8CMRFbsO#C#;R
RRMRC8CRoMNCs0zCR4
6;RRRRzR4n:VRHRF5M0NRI8_8ss2CoRMoCC0sNCR
RRRRRRRRRRNRI8C_so=R<R7Wq7
);RRRRCRM8oCCMsCN0Rnz4;R

R-RR-CRtMNCs00CRE)CRqOvRC#DDR8NMRD#CCRO0DHFoOR
RR4Rz4RR:VRFsHMRHRlMk_DOCD8#RF0IMFRRjoCCMsCN0
RRRRRRRRR--Q5VRNs88I0H8ERR>cM2RCRC80OFRs0CNCsRIHR0CCLMNDNCRMF8Rkk0b0MRCNCLDRD#CCRO0DHFoOR
RRRRRR4Rz.RR:H5VRNs88I0H8ERR>co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4RCIEMsR5Ns8_CNo58I8sHE80-84RF0IMF2RcRH=R2DRC#'CRj
';RRRRRRRRRRRRRRRRI_s0CHM52=R<RRW IMECRN5I8C_so85N8HsI8-0E4FR8IFM0RRc2=2RHR#CDCjR''R;
RRRRRCRRMo8RCsMCNR0Cz;4.
RRRRRRRRR--Q5VRNs88I0H8E=R<RRc2MIFRsCH0RNCMLRDCFFsRkk0b0MRCNCLDRD#CCRO0DHFoOCRMC88C
RRRRRRRRdz4RH:RVNR58I8sHE80RR<=co2RCsMCN
0CRRRRRRRRRRRRRRRRF_k0CHM52=R<R''4;R
RRRRRRRRRRRRRRsRI0M_C5RH2<W=R R;
RRRRRRRRRCRRMo8RCsMCNR0Cz;4d
RRRRR--tsMCNR0C0REC)RqvODCD#MRN8sR0H0-#N#0C
RRRRRRRRcz4RV:RF[sRRRHM58IH0-ERRR428MFI0jFRRMoCC0sNCR
RRRRRRRRRR0RN0LsHkR0C\N3slV_FV0#C\VRFRqz)vRR:DCNLD#RHR7"1a&"RR0HMCsoC'NHloIC5HE802RR&"R7"&MRH0CCosl'HN5oCHn*42RR&"RW"&MRH0CCosl'HN5oC[&2RR"" RH&RMo0CCHs'lCNo50oC_8CM_b8C05E5H2+4*,4nRb8C02E2R"&RX&"RR0HMCsoC'NHlo[C5+;42
RRRRRRRRRRRRoLCHRM
RRRRRRRRRzRR):qvRv)q44nX7RR
RRRRRRRRRRRRRbRRFRs0lRNb5=7R>MRH_osC5,[2RRqj=D>RFII_Ns885,j2RRq4=D>RFII_Ns885,42RRq.=D>RFII_Ns885,.2
RRRRRRRRRRRRRRRRRRRRRRRRqRRd>R=RIDF_8IN8ds527,Ruj)qRR=>D_FIs8N8s25j,uR7)Rq4=D>RFsI_Ns885,42RR
RRRRRRRRRRRRRRRRRRRRRRRRR7qu).>R=RIDF_8sN8.s527,Rud)qRR=>D_FIs8N8s25d, RWRR=>I_s0CHM52
,RRRRRRRRRRRRRRRRRRRRRRRRRRBRWp=iR>pRBi7,Ru=mR>kRF0k_L#,5H[;22
RRRRRRRRRRRR0Fk_osC5R[2<F=RkL0_kH#5,R[2IMECRk5F0M_C5RH2=4R''C2RDR#C';Z'
RRRRRRRRRRRR8CMRMoCC0sNC4RzcR;
RRRRRCRRMo8RCsMCNR0Cz;44
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR
MN8RsHOE00COkRsC#CCDOs0_N
l;
