@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
`RRHDMOkR8C"8#0_DFP_#0N	"3E
R
RbNNslCC0s#RN#0Cs_lMNCRR="1q1 _)aQ)hB hv a
";
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_BQh)  vhua_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5#L0ND0C5C_#0CsGb2&2R&bRfN5#0`pme_1)  1a_Qqthp22RR>|-R55R00C#_bCGsRR>f#bN0C50#C0_G2bs2
R?RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RR00C#_bCGsRR-f#bN0C50#C0_G2bsRR==PkNDC:2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5#0C0G_Cb+sRRI5{HE80{L4'4R}}-bRfN5#000C#_bCGsR22+'R4L=4R=NRPD2kC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2R;
R8CMbbsFC$s0
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRsRbFsbC0q$R1)1 ah_QBv)  _haXmZ_h _a1 a_X_u)uR;
RR@@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R!R55#fHkMM	F5IM00C#_bCGs222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
CR
RRRR#ONCbR5sCFbs_0$0C$b2R
RRRRR`pme_1q1 R)a:CRLoRHM:PRFD#_N#0Cs
RRRRRRRRqq_1)1 ah_QBv)  _hauR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )_BQh)  vhua_2DRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMHH#RMCOsN8#CRRL$NNRPDRkCFC0EsER0N#MRbHCOV8HC"
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)Qa_h B)va h__XZmah_ _1a )Xu_
u:RRRRRRRRNC##sb0RsCFbsR0$51q1 _)aQ)hB hv aZ_X__mhaa 1_u X)2_u
RRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R

RRRRRe`mp1_q1 zvRL:RCMoHRF:RPND_#l#kCR
RRRRRR_Rvq 11)Qa_h B)va h_Ru:Nk##lbCRsCFbsR0$51q1 _)aQ)hB hv a2_u;
R
`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqv_1)1 ah_QBv)  _haXmZ_h _a1 a_X_u)uR:
RRRRRNRR#l#kCsRbFsbC05$Rq 11)Qa_h B)va h__XZmah_ _1a )Xu_;u2
`RRCHM8V/R/m_epQpvuQaBQ_]XB _Bim
ww`8CMH/VR/pme_]XB _Bim
ww
RRRRCRRMR8
RRRRRe`mpt_Qh m)RL:RCMoHRF:RPHD_osMFCR
RRRRRR/R/RR8FMEF0HRMo;R
RRRRRC
M8RRRRRCR8VDNk0RRRRRR:H0MHHRNDF_PDCFsss5_0";"2
RRRR8CMOCN#
R
RCoM8CsMCN
0C
M`C8RHV/m/Reqp_1)1 ah_m
H
`VV8CRpme_eBm m)_hR

RMoCC0sNCR

RHRRVOR5FsPCN_oCDCCPD=R!Re`mpm_Be_ )h mh2CRLoRHM:PRFDF_OP
CsRRRRRRHV5pme_eBm A)_qB1Q_2mhRoLCH:MRRDFP_POFCLs_NO#H
R
RRRRROCFPsC_0#C0_G_bsOMENo
C:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRfR!#L0ND0C5C_#0CsGb22R2
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_NOEMRoCOCFPs"C82R;
RRRRC
M8RRRRC
M8
CRRMC8oMNCs0
C
`8CMH/VR/eRmpm_Be_ )m
h

