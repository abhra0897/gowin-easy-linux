@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ha_m)_aqQh1ahQm"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
H
`VV8CRpme_QQha1_vtR
RRMRHHN0HDR
RRRRRF_PDH0MH_ol#_R0;/B/RNRDD0RECzs#CRV7CH8MCRHQM0CRv#o#NCFR)kM0HCC
`MV8HRm//eQp_h_Qav
1t
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )__hmah)q1QQamuh_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5#0C0G_Cb=sR=0R#N_s0#00NC|2R=5>R00C#_bCGs=R!RNfb#M05C_G0#00NC;22
CRRMs8bFsbC0
$

V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RbbsFC$s0R1q1 _)aham_)1qhQmaQhZ_X__mhaa 1_u X);_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR55!fkH#MF	MI0M5C_#0CsGb2;22
CRRMs8bFsbC0
$
RsRbFsbC0q$R1)1 am_h_qa)ha1QQ_mhXmZ_ha_1q_)a1aaq ;_u
@RR@F5b#oC8CDRO	R2
R#8HNCLDRVHVRm5`e)p_ a1 _t1QhRqp!4=R'2L4
RRRR55!fkH#MF	MI#M500Ns_N#002C22R;
R8CMbbsFC$s0
R
RbbsFC$s0R1q1 _)aham_)1qhQmaQhZ_X__mhha X_q1aau _;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
RR0R5C_#0CsGbRR==#s0N00_#N20CR>|-R55!fkH#MF	MIMM5C_G0#00NC222;R
RCbM8sCFbs
0$RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RCRoMNCs0
C
RRRROCN#Rs5bFsbC00$_$2bC
RRRR`RRm_epq 11):aRRoLCH:MRRDFP_#N#C
s0RRRRRRRRq1_q1a )__hmah)q1QQamuh_:#RN#0CsRFbsb0Cs$qR51)1 am_h_qa)ha1QQ_mhuR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCPRFDs_Cs_Fs0a5"CR#0CsGbCH##F0MRs#NMHF0HMRC8VlsFRDPNkCCRJDkNRR0F#s0N00_#NR0C0NFRRDPNkCCRJDkNRR0FM0CG_N#002C";


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
RRRRRRRRqq_1)1 am_h_qa)ha1QQ_mhXmZ_h _a1 a_X_u)uR:
RRRRRRRRR#N#CRs0bbsFC$s0R15q1a )__hmah)q1QQamXh_Zh_m_1a aX_ uu)_2R
RRRRRRRRRCCD#RDFP_sCsF0s_5C"0#C0_GRbsO0FMN#HMRFXRs"RZ2
;
RRRRRRRRq1_q1a )__hmah)q1QQamXh_Zh_m_q1a)1a_a qa_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 am_h_qa)ha1QQ_mhXmZ_ha_1q_)a1aaq 2_u
RRRRRRRRCRRDR#CF_PDCFsss5_0"N#0s#0_0CN0RMOF0MNH#RRXFZsR"
2;
RRRRRRRRqq_1)1 am_h_qa)ha1QQ_mhXmZ_h _hX1a_a qa_
u:RRRRRRRRR#RN#0CsRFbsb0Cs$qR51)1 am_h_qa)ha1QQ_mhXmZ_h _hX1a_a qa_
u2RRRRRRRRRDRC#FCRPCD_sssF_"05M0CG_N#00OCRFNM0HRM#XsRFR2Z";R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw



RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRqv_1)1 am_h_qa)ha1QQ_mhuN:R#l#kCsRbFsbC05$Rq 11)ha_m)_aqQh1ahQm_;u2
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )__hmah)q1QQamXh_Zh_m_1a aX_ uu)_:R
RRRRRRRRRNk##lbCRsCFbsR0$51q1 _)aham_)1qhQmaQhZ_X__mhaa 1_u X)2_u;R

RRRRRvRR_1q1 _)aham_)1qhQmaQhZ_X__mh1)aqaa_1q_a uR:
RRRRRRRRR#N#kRlCbbsFC$s0R15q1a )__hmah)q1QQamXh_Zh_m_q1a)1a_a qa_;u2
R
RRRRRR_Rvq 11)ha_m)_aqQh1ahQm__XZmhh_ _Xa1aaq :_u
RRRRRRRRNRR#l#kCsRbFsbC05$Rq 11)ha_m)_aqQh1ahQm__XZmhh_ _Xa1aaq 2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw



RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//8MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
V`H8RCVm_epB me)h_m
C
oMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR

RRRRRPOFC#s_00Ns_N#00
C:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRR5#0C0G_Cb=sR=0R#N_s0#00NCR222R
RRRRRRRRRRRRRRRRRRFRRPOD_FsPC_"05#s0N00_#NR0COCFPs"C82R;
RRRRC
M8RRRRC
M8
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m
