@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)Wa_Q]7a"
;
RHR`MkOD8"CR#_08F_PD0	N#3
E"
V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
RMRHHN0HDCRLo
HMRRRRH5VRRH5lM	_O#RR>j&2R&lR5NOG_	>#RRRj22CRLo
HMRRRRRVRHRH5lM	_O#RR>l_NGO2	#RDFP_sCsF0s_5D"QDNCoDNRbsCNl0RCsPkNDC##RCI0RECCsRMlH_#O	Rl>RNOG_	2#";R
RRMRC8R
RC
M8
V`H8RCVm_epq 11)ma_hR

RFbsb0Cs$1Rq1a )_7WQav]_QBh_]i B_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42RsRfF5#C00C#_bCGs|2R-5>R00C#_bCGslr*HOM_	2#9;R
RCbM8sCFbs
0$
bRRsCFbsR0$q 11)Wa_Q]7a_Xvq_ B]Bui_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
Rf#sFCC50#C0_G2bsR>|-RC50#C0_Grbs*54:l_NGOR	#>RRj?NRlG	_O#RR:.229R4yyR05!C_#0CsGb2R;
R8CMbbsFC$s0
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RFbsb0Cs$1Rq1a )_7WQaX]_Zh_m_1a aX_ uu)_;R
R@b@5F8#CoOCRD
	2RHR8#DNLCVRHV`R5m_ep)  1aQ_1tphqRR!=44'L2R
R5f!5HM#k	IMFMC50#C0_G2bs2
2;RMRC8Fbsb0Cs$R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RoCCMsCN0
R
RRNRO#5CRbbsFC$s0_b0$CR2
RRRRRe`mp1_q1a )RL:RCMoHRF:RPND_#s#C0R
RRRRRRVRHRH5lM	_O#RR>jL2RCMoHRN:R_#N#C_s0I0H8EH_lME_OC
O	RRRRRRRRR_Rqq 11)Wa_Q]7a_hvQ_ B]Bui_:#RN#0CsRFbsb0Cs$qR51)1 aQ_W7_a]v_QhBB] i2_u
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRDR#CF_PDCFsss5_0"#aC0GRCb#sC#MHFR#INRDEC8)RazV RFDsRCR##0MENRC#bOHHVCl8RHlMHkllRHOM_	O#R$COD#;"2
RRRRRRRR8CM
RRRRRRRRRHV5GlN_#O	Rj>R2CRLoRHM:_RNNC##sI0_HE80_GlN_COEOR	
RRRRRRRRRqq_1)1 aQ_W7_a]v_qXBB] i:_uR#N#CRs0bbsFC$s0R15q1a )_7WQav]_qBX_]i B_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRDRC#FCRPCD_sssF_"05a0C#RbCGs#C#HRFMIRN#E8CDRza) FRVsFRls0CRERNM#ObCHCVH8NRlGkHllNRlG	_O#$ROO#DC"
2;RRRRRRRRC
M8
H
`VV8CRpme_]XB _Bim
wwR/R/7MFRFH0EM`o
CCD#
`RRHCV8VeRmpv_QuBpQQXa_BB] iw_mwR
RR/R/7MFRFH0EMRo
RD`C#RC
RRRRRRRRq1_q1a )_7WQaX]_Zh_m_1a aX_ uu)_:R
RRRRRRNRR#s#C0sRbFsbC05$Rq 11)Wa_Q]7a__XZmah_ _1a )Xu_
u2RRRRRRRRR#CDCPRFDs_Cs_Fs005"C_#0CsGbRMOF0MNH#RRXFZsR"
2;RCR`MV8HRm//eQp_vQupB_QaX B]Bmi_w`w
CHM8V/R/m_epX B]Bmi_w
w
RRRRRMRC8R
RRRRR`pme_1q1zRv :CRLoRHM:PRFD#_N#Ckl
RRRRRRRRRHV5MlH_#O	Rj>R2CRLoRHM:_RlNC##sI0_HE80_MlH_COEOR	
RRRRRRRRRqv_1)1 aQ_W7_a]v_QhBB] i:_uR#N#kRlCbbsFC$s0R15q1a )_7WQav]_QBh_]i B_;u2
RRRRRRRR8CM
RRRRRRRRRHV5GlN_#O	Rj>R2CRLoRHM:_RlNC##sI0_HE80_GlN_COEOR	
RRRRRRRRRqv_1)1 aQ_W7_a]v_qXBB] i:_uR#N#kRlCbbsFC$s0R15q1a )_7WQav]_qBX_]i B_;u2
RRRRRRRR8CM
`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRRqv_1)1 aQ_W7_a]XmZ_h _a1 a_X_u)uR:
RRRRRRRRNk##lbCRsCFbsR0$51q1 _)aWaQ7]Z_X__mhaa 1_u X)2_u;R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R
RRRRRC
M8RRRRRmR`eQp_t)hm RR:LHCoMRR:F_PDHFoMsRC
RRRRR/RR/FR8R0MFEoHMRR;
RRRRR8CM
RRRR8RRCkVNDR0RR:RRRHHM0DHNRDFP_sCsF0s_52"";R
RRMRC8#ONCR

R8CMoCCMsCN0
C
`MV8HRR//m_epq 11)ma_h`

HCV8VeRmpm_Be_ )m
h
oCCMsCN0
R
RRVRHRF5OPNCsoDC_CDPCRR!=`pme_eBm h)_m2h RoLCH:MRRDFP_POFCRs
RRRRH5VRm_epB me)q_A1_QBmRh2LHCoMRR:F_PDOCFPsN_L#
HO
RRRRORRFsPC_#0C0G_CbNs_#s#C0
#:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRfF5#C00C#_bCGsR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2R
RRRRRRRRRRRRRRRRRR2RR
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_#N#C#s0RPOFC8sC"
2;RRRRR8CM
R
RRHRRVmR5eBp_m)e _)Bmh_ )mRh2LHCoMRR:F_PDOCFPsF_OssMC
RRRRHRRVlR5HOM_	>#RRRj2LHCoMRR:F_PDOCFPsC_0#C0_G_bsNC##s80C_sVF_MlH_#O	
RRRRRRR
RRRRRRROCFPsC_0#C0_G_bsNC##s80C_sVF_MlH_#O	:R
RRRRRRPOFCbsRsCFbsR0$55@@bCF#8RoCO2D	Rm5`e)p_ a1 _t1QhRqp!4=R'2LjRs0EFEkoF
k0RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRfR5sCF#5#0C0G_Cb
s2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRyRyjR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5#0C0G_Cb*srl_HMO9	#2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRy
y4RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR!R500C#_bCGsR2
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR2R
RRRRRRRRRRRRRRRRRRRRR2R
RRRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbNs_#s#C0_C8V_Fsl_HMOR	#OCFPs"C82R;
RRRRR8CM
R
RRRRRH5VRl_NGOR	#>2RjRoLCH:MRRDFP_POFC0s_C_#0CsGb_#N#CCs08F_VsN_lG	_O#R
RRRR
RRRRRFROP_Cs00C#_bCGs#_N#0CsCV8_Fls_NOG_	
#:RRRRRORRFsPCRFbsb0Cs$@R5@F5b#oC8CDRO	52R`pme_1)  1a_Qqthp=R!RL4'j02REksFokEF0R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5Ffs#0C5C_#0CsGb2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRy
yjRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0R5C_#0CsGbrN*lG	_O#
92RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRyRy4R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5C!0#C0_G2bs
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR
R2RRRRRRRRRRRRRRRRRRRRR
R2RRRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb_#N#CCs08F_VsN_lG	_O#FROPCCs8;"2
RRRRCRRM
8
RRRRR8CMRO//FCsMsFROPNCsoRC
RCRRM
8
CoM8CsMCN
0C
M`C8RHV/m/ReBp_m)e _
mh
