`ifndef ATCAPBBRG100_CONST_VH
`define ATCAPBBRG100_CONST_VH

`include "ae250_config.vh"
`include "ae250_const.vh"

`define	ATCAPBBRG100_PRODUCT_ID			32'h00021008

`ifdef ATCAPBBRG100_ADDR_WIDTH_24
`define	ATCAPBBRG100_ADDR_MSB			23
`define ATCAPBBRG100_SLV_OFFSET_UNIT		10
`else
`define	ATCAPBBRG100_ADDR_MSB			31
`define ATCAPBBRG100_SLV_OFFSET_UNIT		20
`endif

`define ATCAPBBRG100_SPACE_MSB			(`ATCAPBBRG100_ADDR_DECODE_WIDTH - 1)

`define ATCAPBBRG100_SLV_0

`ifdef ATCAPBBRG100_ADDR_WIDTH_24
`define ATCAPBBRG100_SLV0_SIZE			3
`else
`define ATCAPBBRG100_SLV0_SIZE			1
`endif

`ifndef ATCAPBBRG100_SLV0_OFFSET
`define	ATCAPBBRG100_SLV0_OFFSET		`ATCAPBBRG100_ADDR_DECODE_WIDTH'h0
`endif

`define ATCAPBBRG100_SLV0_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV0_SIZE - 1)
`define ATCAPBBRG100_SLV1_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV1_SIZE - 1)
`define ATCAPBBRG100_SLV2_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV2_SIZE - 1)
`define ATCAPBBRG100_SLV3_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV3_SIZE - 1)
`define ATCAPBBRG100_SLV4_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV4_SIZE - 1)
`define ATCAPBBRG100_SLV5_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV5_SIZE - 1)
`define ATCAPBBRG100_SLV6_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV6_SIZE - 1)
`define ATCAPBBRG100_SLV7_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV7_SIZE - 1)
`define ATCAPBBRG100_SLV8_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV8_SIZE - 1)
`define ATCAPBBRG100_SLV9_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV9_SIZE - 1)
`define ATCAPBBRG100_SLV10_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV10_SIZE - 1)
`define ATCAPBBRG100_SLV11_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV11_SIZE - 1)
`define ATCAPBBRG100_SLV12_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV12_SIZE - 1)
`define ATCAPBBRG100_SLV13_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV13_SIZE - 1)
`define ATCAPBBRG100_SLV14_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV14_SIZE - 1)
`define ATCAPBBRG100_SLV15_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV15_SIZE - 1)
`define ATCAPBBRG100_SLV16_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV16_SIZE - 1)
`define ATCAPBBRG100_SLV17_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV17_SIZE - 1)
`define ATCAPBBRG100_SLV18_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV18_SIZE - 1)
`define ATCAPBBRG100_SLV19_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV19_SIZE - 1)
`define ATCAPBBRG100_SLV20_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV20_SIZE - 1)
`define ATCAPBBRG100_SLV21_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV21_SIZE - 1)
`define ATCAPBBRG100_SLV22_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV22_SIZE - 1)
`define ATCAPBBRG100_SLV23_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV23_SIZE - 1)
`define ATCAPBBRG100_SLV24_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV24_SIZE - 1)
`define ATCAPBBRG100_SLV25_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV25_SIZE - 1)
`define ATCAPBBRG100_SLV26_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV26_SIZE - 1)
`define ATCAPBBRG100_SLV27_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV27_SIZE - 1)
`define ATCAPBBRG100_SLV28_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV28_SIZE - 1)
`define ATCAPBBRG100_SLV29_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV29_SIZE - 1)
`define ATCAPBBRG100_SLV30_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV30_SIZE - 1)
`define ATCAPBBRG100_SLV31_OFFSET_LSB		(`ATCAPBBRG100_SLV_OFFSET_UNIT + `ATCAPBBRG100_SLV31_SIZE - 1)
`define ATCAPBBRG100_OFFSET_MSB			`ATCAPBBRG100_SPACE_MSB


`define ATCAPBBRG100_SLV1_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV1_OFFSET} | 33'd`ATCAPBBRG100_SLV1_SIZE)
`define ATCAPBBRG100_SLV2_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV2_OFFSET} | 33'd`ATCAPBBRG100_SLV2_SIZE)
`define ATCAPBBRG100_SLV3_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV3_OFFSET} | 33'd`ATCAPBBRG100_SLV3_SIZE)
`define ATCAPBBRG100_SLV4_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV4_OFFSET} | 33'd`ATCAPBBRG100_SLV4_SIZE)
`define ATCAPBBRG100_SLV5_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV5_OFFSET} | 33'd`ATCAPBBRG100_SLV5_SIZE)
`define ATCAPBBRG100_SLV6_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV6_OFFSET} | 33'd`ATCAPBBRG100_SLV6_SIZE)
`define ATCAPBBRG100_SLV7_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV7_OFFSET} | 33'd`ATCAPBBRG100_SLV7_SIZE)
`define ATCAPBBRG100_SLV8_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV8_OFFSET} | 33'd`ATCAPBBRG100_SLV8_SIZE)
`define ATCAPBBRG100_SLV9_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV9_OFFSET} | 33'd`ATCAPBBRG100_SLV9_SIZE)
`define ATCAPBBRG100_SLV10_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV10_OFFSET} | 33'd`ATCAPBBRG100_SLV10_SIZE)
`define ATCAPBBRG100_SLV11_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV11_OFFSET} | 33'd`ATCAPBBRG100_SLV11_SIZE)
`define ATCAPBBRG100_SLV12_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV12_OFFSET} | 33'd`ATCAPBBRG100_SLV12_SIZE)
`define ATCAPBBRG100_SLV13_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV13_OFFSET} | 33'd`ATCAPBBRG100_SLV13_SIZE)
`define ATCAPBBRG100_SLV14_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV14_OFFSET} | 33'd`ATCAPBBRG100_SLV14_SIZE)
`define ATCAPBBRG100_SLV15_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV15_OFFSET} | 33'd`ATCAPBBRG100_SLV15_SIZE)
`define ATCAPBBRG100_SLV16_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV16_OFFSET} | 33'd`ATCAPBBRG100_SLV16_SIZE)
`define ATCAPBBRG100_SLV17_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV17_OFFSET} | 33'd`ATCAPBBRG100_SLV17_SIZE)
`define ATCAPBBRG100_SLV18_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV18_OFFSET} | 33'd`ATCAPBBRG100_SLV18_SIZE)
`define ATCAPBBRG100_SLV19_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV19_OFFSET} | 33'd`ATCAPBBRG100_SLV19_SIZE)
`define ATCAPBBRG100_SLV20_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV20_OFFSET} | 33'd`ATCAPBBRG100_SLV20_SIZE)
`define ATCAPBBRG100_SLV21_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV21_OFFSET} | 33'd`ATCAPBBRG100_SLV21_SIZE)
`define ATCAPBBRG100_SLV22_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV22_OFFSET} | 33'd`ATCAPBBRG100_SLV22_SIZE)
`define ATCAPBBRG100_SLV23_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV23_OFFSET} | 33'd`ATCAPBBRG100_SLV23_SIZE)
`define ATCAPBBRG100_SLV24_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV24_OFFSET} | 33'd`ATCAPBBRG100_SLV24_SIZE)
`define ATCAPBBRG100_SLV25_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV25_OFFSET} | 33'd`ATCAPBBRG100_SLV25_SIZE)
`define ATCAPBBRG100_SLV26_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV26_OFFSET} | 33'd`ATCAPBBRG100_SLV26_SIZE)
`define ATCAPBBRG100_SLV27_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV27_OFFSET} | 33'd`ATCAPBBRG100_SLV27_SIZE)
`define ATCAPBBRG100_SLV28_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV28_OFFSET} | 33'd`ATCAPBBRG100_SLV28_SIZE)
`define ATCAPBBRG100_SLV29_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV29_OFFSET} | 33'd`ATCAPBBRG100_SLV29_SIZE)
`define ATCAPBBRG100_SLV30_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV30_OFFSET} | 33'd`ATCAPBBRG100_SLV30_SIZE)
`define ATCAPBBRG100_SLV31_CFG_REG		({{33-`ATCAPBBRG100_ADDR_DECODE_WIDTH{1'b0}}, `ATCAPBBRG100_SLV31_OFFSET} | 33'd`ATCAPBBRG100_SLV31_SIZE)
`define ATCAPBBRG100_REG_ADDR_WIDTH		8
`define	ATCAPBBRG100_REG_ADDR_MSB		(`ATCAPBBRG100_REG_ADDR_WIDTH + 1)

`endif
