@ER//qCOODsDCN0R1NNM8se8R4R3UmMbCRseCHOVHNF0HMHRpLssN$mR5e3p2
R//qCOODsDCNFRBbH$soRE05RO2.6jj-j.jnq3RDsDRH0oE#CRs#PCsC
83
bRRNlsNCs0CR#N#C_s0MCNlR"=Rq 11)ha_mh_z7w )p"mW;R

RM`HO8DkC#R"0F8_P0D_N3#	E
"

V`H8RCVm_epQahQ_tv1
RRRRHHM0DHN
RRRRFRRPHD_M_H0l_#o0/;R/NRBD0DREzCR#RCs7HCVMRC8Q0MHR#vC#CNoRk)F0CHM
M`C8RHV/e/mph_QQva_1
t
`8HVCmVReqp_1)1 ah_m
R
RbbsFC$s0R1q1 _)ahzm_h)7 wWpm_
u;R@R@5#bFCC8oR	OD2R
R8NH#LRDCHRVV5e`mp _)1_ a1hQtq!pR='R4L
42R0R5C_#0CsGbRR==l2HMR>|=R055C_#0CsGbRl<RNRG2&5&R00C#_bCGs=R>RMlH2
2;RMRC8Fbsb0Cs$


`8HVCmVReXp_BB] iw_mwR
R/F/7R0MFEoHM
D`C#RC
RV`H8RCVm_epQpvuQaBQ_]XB _Bim
wwRRRR/F/7R0MFEoHM
`RRCCD#
bRRsCFbsR0$q 11)ha_mh_z7w )p_mWXmZ_h _a1 a_X_u)uR;
R5@@bCF#8RoCO2D	
8RRHL#NDHCRV5VR`pme_1)  1a_Qqthp=R!RL4'4R2
R55!fkH#MF	MI0M5C_#0CsGb2;22
CRRMs8bFsbC0R$
RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mwR

RMoCC0sNCR

RORRNR#C5Fbsb0Cs$$_0b
C2RRRRRmR`eqp_1)1 aRR:LHCoMRR:F_PDNC##sR0
RRRRRqRR_1q1 _)ahzm_h)7 wWpm_Ru:NC##sb0RsCFbsR0$51q1 _)ahzm_h)7 wWpm_
u2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#CDCPRFDs_Cs_Fs0a5"CR#0CsGbCH##FOMREoNMCP8RNCDkRFVslDRNDCFI8HRlMkHllNRPDRkClRHM0NFRRDPNkHCRMER0CNRsMRoCl-HM4FR0RGlN"
2;
V`H8RCVm_epX B]Bmi_wRw
R7//FFRM0MEHoC
`D
#CRHR`VV8CRpme_uQvpQQBaB_X]i B_wmw
RRRR7//FFRM0MEHoR
R`#CDCR
RRRRRR_Rqq 11)ha_mh_z7w )p_mWXmZ_h _a1 a_X_u)uR:
RRRRRNRR#s#C0sRbFsbC05$Rq 11)ha_mh_z7w )p_mWXmZ_h _a1 a_X_u)uR2
RRRRRCRRDR#CF_PDCFsss5_0"#0C0G_CbOsRFNM0HRM#XsRFR2Z";R
R`8CMH/VR/pme_uQvpQQBaB_X]i B_wmw
M`C8RHV/e/mpB_X]i B_wmw
R

RRRRR8CM
RRRR`RRm_epqz11v: RRoLCH:MRRDFP_#N#k
lCRRRRRRRRv1_q1a )__hmz h7)mwpW:_uR#N#kRlCbbsFC$s0R15q1a )__hmz h7)mwpW2_u;`

HCV8VeRmpB_X]i B_wmw
/RR/R7FMEF0H
Mo`#CDCR
R`8HVCmVReQp_vQupB_QaX B]Bmi_wRw
R/RR/R7FMEF0H
MoRCR`D
#CRRRRRRRRv1_q1a )__hmz h7)mwpWZ_X__mhaa 1_u X):_u
RRRRRRRR#N#kRlCbbsFC$s0R15q1a )__hmz h7)mwpWZ_X__mhaa 1_u X)2_u;R

RM`C8RHV/e/mpv_QuBpQQXa_BB] iw_mwC
`MV8HRm//eXp_BB] iw_mw


RRRRRMRC8R
RRRRR`pme_hQtmR) :CRLoRHM:PRFDo_HMCFs
RRRRRRRRR//7MFRFH0EM;oR
RRRRCRRMR8
RRRRRV8CN0kDRRRRRH:RMHH0NFDRPCD_sssF_"05"
2;RRRRCOM8N
#C
CRRMC8oMNCs0
C
`8CMH/VR/eRmp1_q1a )_
mh
V`H8RCVm_epB me)h_m
C
oMNCs0
C
RRRRH5VROCFPsCNo_PDCC!DR=mR`eBp_m)e _hhm L2RCMoHRF:RPOD_FsPC
RRRRVRHRe5mpm_Be_ )AQq1Bh_m2CRLoRHM:PRFDF_OP_CsLHN#OR
RR
RRRRRRRFROP_Cs00C#_bCGs0_N_MlH:R
RRRRROCFPssRbFsbC05$R@b@5F8#CoOCRDR	25`R5m_ep)  1aQ_1tphqRR!=4j'L2&R&
RRRRRRRRRRRRRRRRRRRRsRfF5#C00C#_bCGs=R=RMlH22R2
RRRRRRRRRRRRRRRRRRRRPRFDF_OP_Cs005"C_#0CsGb__N0lRHMOCFPs"C82R;
RRRRCRM8/N/L#RHOOCFPsCCo
R
RRHRRVmR5eBp_m)e _)Bmh_ )mRh2LHCoMRR:F_PDOCFPsF_OssMC
R
RRRRROCFPsC_0#C0_G_bsNl0_N
G:RRRRRFROPRCsbbsFC$s0R@5@5#bFCC8oR	OD2RR55e`mp _)1_ a1hQtq!pR='R4LRj2&R&
RRRRRRRRRRRRRRRRRRRRf#sFCC50#C0_GRbs=l=RNRG22R2
RRRRRRRRRRRRRRRRRRRRF_PDOCFPs5_0"#0C0G_CbNs_0N_lGFROPCCs8;"2
RRRRMRC8/R/OMFsCOsRFsPCN
oCRRRRC
M8
8CMoCCMsCN0
C
`MV8HRR//m_epB me)h_m
