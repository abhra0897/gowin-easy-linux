-- This is a customized version of the float_generic_pkg package
@ER--wRFs1b$MD$HVR7e]p$R1MC0E#3H#
-

--R--------------------------------------------------------------------
--
-RbBF$osHE�0RRj.jU$RLR Q  q3RDsDRH0oE#CRs#PCsC
83---
-ERaH##RFOksCHRVDHCR#MRNR#C#CHM0NbDRNRs0FQVR R  1R084nj(-j.jU-,
- RQ 1 R08NMNRs8ep]7RMpNookNCCR)VCCsMROCvkNMNRD3a#EHRk#FsROCVCHDR$lNR0MFR
LC-O-RFCbH8#,RF,D8RRFsHDMOk88CR0IHEFR#VN0Is0CRERN0H##RFRD8IEH0FRk0I0sH0RCM
R--blCsHH##FVMRsRFl0RECQ   RN10Ms8N87#RCsbN0MlC0a3RERH##sFkOVCRHRDClRN$L
CR-O-RFCbH8FRVsMRH8HHP8DkNRCk#R0LCIMCCRODHCCM#8#RkC3s#RHaE#FR#kCsORDVHC#RH
R--bPsFH88CRRFMNqMR11RQR#LNHR#3aRECQ   R#8HOHDNlq#RhWYRqq))hRaY )Xu R11m-)
-vRQu pQ7hRQB7pzQRhtqRhYW)q)qYhaRRmwvB )]aqhqpAQQRaYqRh7whQa R11wRm)z
1 -w-Rmq)RR)uqazQBpRq)uuz)m31 RCaERCk#sVRFRC0ERk#FsROCVCHDRN#EDHDRMl8CM$HV
R--NRM8E8FDR Q  NREsClD#V#RsRFlNRM$8NNloRC#FDsRHHNLD$H0RHNs#oHMR0FkRRFV0
EC-k-R#0CRECCsF
V3---
-RRRaDH0CRRRRRR:RFwDNM0HoF-bHRM0b	NONRoC5MtCCOsHRObN	CNoRO8CDNNs0MHF2-
-RRRRRRRRRRRRR-:
-RRRpsHLNRs$RRR:RHaE#NRbOo	NCER#NRDDLOCRFHlbDRC8HFM0RDNRHNLss-$
-RRRRRRRRRRRRRR:Rl#$LHFDODND$NRMlRC8Q   3-
-RRRRRRRRRRRRR-:
-RRR7CCPDCFbsR#:ROqOCCDDseNR]-7paNBRMQ8R R  u(4jnFRWsM	HosRtF
kb-R-RRRRRRRRRR:RR
R--RkRus#bFCRRR:aRRERH#b	NON#oCRV8CH#MCR#LNHLORHsMN$DRVFHN0MboRF0HM
R--RRRRRRRRRRRR:NRRsEH0lHC0OkRVMHO0F
M#-R-RRRRRRRRRR:RR
R--RFRh0RCRRRRR:aRRERH#b	NONRoClRN$LlCRFV8HHRC80HFRMkOD8NCR808HHNFMDNR80-N
-RRRRRRRRRRRRRR:RJsCkCHs8$RLRF0FDR#,LRk0Hl0RkR#0HMMRFNRI$ERONCMoRC0E
R--RRRRRRRRRRRR:CRRGs0CMRNDHCM0sOVNCF#RsHR#lNkD0MHFRELCNFPHsVRFRC0E
R--RRRRRRRRRRRR:8RRCs#OHHb0FRM3QH0R#CRbs#lH#DHLCFR0R8N8RlOFl0CM#MRN8s/F
R--RRRRRRRRRRRR:NRR0H0sLCk0#FR0RC0ERObN	CNoRO8CDNNs0MHF#L,RkM0RF00RFERONCMo
R--RRRRRRRRRRRR:FRRsCR8DCC0R$NMRHFsoNHMDHRDMRC#F0VREbCRNNO	o8CRCNODsHN0F
M3-R-RRRRRRRRRR:RRRERaCNRbOo	NCFRL8l$RNL$RCERONCMo8MRFDH$RMORNO8FsNCMOR0IHE-
-RRRRRRRRRRRRRR:R0REC0lCs#VRFRNBDkR#C4FnRVER0H##R08NMN3s8
R--RRRRRRRRRRRR:-
-R---------------------------------------------------------------------
-RCf)PHH#FRM:4j..R-f
-7RfN:0CRj.jUc-j-R4j44(:ng:jRg+jd5jRa,EkRR4jqRbs.Ujj2
Rf---R-----------------------------------------------------------------
--
Ck#R71a3Xa a3QmN;DD
LDHs$NsR Q  k;
#QCR 3  1_a7pQmtB4_4nNc3D
D;kR#CQ   3vhz B)Q_71a3DND;#
kC RQ V 3H8GC_FVDN00_$#bC3DND;#
kCCRHCVC3H8GC_ob	3DND;b

NNO	oVCRD0FN_MoCCOsH_ob	R
H#RCRoMHCsO
R5RRRR-7-RCkVNDR0#VRFs#HHxMsoRFHk0M,C#RCIEMFR$kFR8R"NR0VF_D0FN"ER0HI#RHRDDLRC
R-RR-ER0CCR8VDNk0HR#xRC3RN GlCbDRFVDN.0dRkIFDL8RCRRUNRM8.5dRUFR8IFM0Rd-.2R
RRDRVF_N0CFGbM0CM_8IH0:ERRahqzp)qRRRR:U=R;R
RRDRVF_N0VOsN0MHF_8IH0:ERRahqzp)qRRRR:.=RdR;
R-RR-FR)kHM8MNoRDsoFHl0E,sR"F8kM_NMCs0C#"#RHRV8CN0kD,0RFERCsPHND8NRPD#kC
RRRRR--NRsC"ksFMx8_C"sFRs50kNMO0MHF2",RsMFk8M_HV5"RsMFk8bRk2N,RMR8
R-RR-sR"F8kM_oMCH"MVRF5skRM88MFI2R
RRDRVF_N0sMFk80_#$RDCR:RRRksFM08_$RbC:s=RF8kM_NMCs0C#;R
RR-R-RM7CFNslDkRMlsLC#PR5CRs$#DlNDkRMlsLC#CRMNxsRC2sFRk0sCsRFRDVN#RC
RVRRD0FN_M8CFNslDCHxRRRR:mRAmqp hRRRRR:=0Csk;R
RR-R-RsakMF#RMqRhhsRbF#OC#oHMRM5HPHND8kRMlsLC#MRN8PRFCDsVFRI20CskRRFVV#NDCR
RRDRVF_N0OOEC	s_CsRFsR:RRRmAmph qRRRR:0=Rs;kC
RRRRR--tskN8HRL0N#RsNCR888CRR0F0RECL0F0FFlRVPRCCRs$FsbCNF0HMFRVsFRskHM8M
o3RRRR-N-RMM$RNs0kNMDRkClLsHR5MkOD8oHMRRj2NRsCPHND8R3
RVRRD0FN_NoksL8_HR0#RRRR:qRhaqz)pRRRRR:=dR;
R-RR-VRQRza) 0,RERCM0MksRVFVRsINMoHM#MRFR""XRFbsbNNo0MHF
RRRR_MFIMNsHRMoRRRRRRRRRRR:Apmm RqhR:RR=NRVD
#CR2RR;R

RR--qEk0F7sRN8PHR#AHERFb5H8L#bEF@E@P8FD3s
o2RFROMN#0MB0RF)b$H0oEhHF0O:CRR)1aQRht:R=
R"RRB$FbsEHo0jR.jLUR$ RQ R 3qRDDsEHo0s#RCs#CP3C8"
;
R-R-R0hFCER0N00RERH#H"#RQ hatR )soNMC>R<"0,RERk#H$VRFkkR#NCRR0DHCDsN,ER0C0MRERC
RR--8NCVkRD0soNMCHRIDLDRCQR5hta  D)'F0IRFhRQa  t)F'DIRR+XR2
Rb0$ChRz)m 1p7e _FVDNH0R#sRNsRN$5aQh )t RMsNo<CR>F2RVaR17p_zmBtQ;-RR-NRlH0MR$
bCRDRNHRN#zD_VFRN0Hz#Rh1) m pe7D_VF;N0
R
R#0kL$RbCVNDF0#RHR#sCFCDP8hRz)m 1p7e _FVDN
0;R-R--------------------------------------------------------------------------
--R-R-RCz#RC0ERFVDN00R$RbC08FRCMVHCFR$kFsRIVMRD0FNHRMobMFH0kRMlsLC#R3
RR--asECCkRl#L0RCRRNMNCo0CHPR8HMCFGRsER0CNRbOo	NCI#RHRDDCFssskRF0R3
RR--vHHMlRkl#bkbFCs08#RHRk"#Lb0$CDRVF(N0RRH#VNDF0dR5RI8FMR0F-;d2"R
R-"-R#0kL$RbCVNDF0R4nHV#RD0FNRR5n8MFI0-FRg"2;RRH#bLsFN$LDRC0ERN#lD#DC0R
R-b-Rs0NOHDONRCFMRR0Fk3#C
-RR----------------------------------------------------------------------------
R
R-Q-R R  (R6c#oHMDbCRsHCO#MHF
#RRk$L0bzCRh1) m pe7D_VFdN0.#RHR)zh p1me_ 7VNDF0UR5RI8FMR0F-2.d;R
RNNDH#_RzVNDF0Rd.Hz#Rh1) m pe7D_VFdN0.R;
RL#k0C$bRFVDN.0dRRH#VNDF0UR5RI8FMR0F-2.d;R
R-----------------------------------------------------------------------------R
R-Q-R -  (R6c#oHMDbCRsHCO#MHFRFVDNM0HoFRbH3M0RERaHH#R#RRN"FVDN
0"R-R-RRHMBN,RMN8RRmwpqHaRMFRwsN0sMR3RaRECCFGbM0CMRRH#UHRL0I#RH,8CR8NM
-RR-ER0CsRVNHO0FHMR#dR.R0LH#HRI8RC3RHaE#FRVs0lNRMONRDEF8FRskDoE$RR(8HCOl
NDR-R-Ro8HH30#RMRQVHHM0H$R#*R.*(4.R4=R3d( UMRHRH0E#kRMlsLCR##$03Cl
-RR-ERaCHRL0CRsb#sCCNM00MHFRRH#NV#RFFDDI
#:R-R-Rj4RgnU(6Rcd.g4jU6(nc4d.j(gUnd6c.
4jR-R-R(URnd6c.R4j4c.d6Un(g.j4dnc6(jUg4
.dR-R-RjjRjjjjjRjjjjjjjjjjjjjjjjjjjjjjj
jjR-R-R(URRRRRRRRj-R4RRRRRRRRRRRRRRRRR-
.dR-R-R-+/RCRRGRb3RNVsOF0HMR
R-----------------------------------------------------------------------------R

RR--Q   Rc(6Rk8FLRDCbOsCHF#HMR
R#0kL$RbCz h)1emp V7_D0FNnHcR#hRz)m 1p7e _FVDN50R484RF0IMF6R-.
2;RDRNHRN#zD_VFnN0c#RHR)zh p1me_ 7VNDF0;nc
#RRk$L0bVCRD0FNnHcR#DRVFRN05R448MFI0-FR6;.2
-RR----------------------------------------------------------------------------
-RR- RQ ( -68cRFDkLCsRbC#OHHRFMVNDF0oHMRHbFMR03RHaE##RHR"NR8LFkDVCRD0FN"R
R-H-RM,RBR8NMRwNRpamq*HURMFRwsN0sMR3RaRECCFGbM0CMRRH#4L4RHR0#ICH8,MRN8R
R-0-REVCRs0NOHRFMH6#R.HRL0I#RH38CRERaHV#RFNsl0NROMFREDs8RFEkoD4$R6CR8ONHlDR
R-8-RH0oH#R3RQHMVM$H0RRH#..**jRc(H0MRERH#MLklC#sR$C#0lR3
RR--aRECLRH0ssCbCM#C0HN0FHMR##RNRDVFD#FI:R
R-R-Rd4R.j(gUnd6c.jR4gnU(6.cd4Ujg(cn6dj.4gnU(6.cd4Ujg(cn6dj.4gnU(6.cd4Rj
RR--Rj4RgnU(6.cd44jR.6dcng(Ujd4.c(6nU4gj.6dcng(Ujd4.c(6nU4gj.6dcng(Uj
4.R-R-RRR1         R  wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww
-RR-4R4RR4jRRRRRjRRRR-4RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR6R-.R
R-+-R/R-RCFGbM0CMRRRRVOsN0MHF
-RR----------------------------------------------------------------------------
R
R-Q-R R  UR6c&RRBCCG0M88CRCbsOHH#FRM
RL#k0C$bR)zh p1me_ 7VNDF0U4.RRH#z h)1emp V7_D0FNR654RI8FMR0F-.442R;
RHNDNz#R_FVDN.04U#RHR)zh p1me_ 7VNDF0U4.;R
R#0kL$RbCVNDF0U4.RRH#VNDF04R56FR8IFM0R4-4.
2;R-R--------------------------------------------------------------------------
--R-R-RCaERU4.R0LHRFVDNM0HoFRbHRM0MLklCHsR#DR"FRMo8LFkDRC"HBMRRM5F
-RR-FR#l#CR$C#0l0#RERH#HN#RRR(jLRH0VNDF0oHMRHbFMM0RkClLsN2RMw8Rpamq*
d.R-R-RRHMw0Fss3NMRERaCGRCbCFMMH0R#6R4R0LH#HRI8NCRM08REVCRs0NOHRFMH4#R4R.
RR--L#H0R8IHCa3RERH#MLklCOsRNEMRNDM8CbRNbGsFH0lNCRD$d8dRClOHN8DRH0oH#R3
RR--QHMVM$H0RRH#.d**.n,((MRHRH0E#kRMlsLCR##$03Cl
-RR----------------------------------------------------------------------------
R
R-b-RkFsb#RC:BOEC	V#RFNsRRDPNHV8RD0FNHRMobMFH0kRMlsLC
0RR$RbCPHND8b_V#00NC#RHRN5MMR,RRRRRRRRRRR--1MHoNMDHoNRhhBR5R_wuh2qh
RRRRRRRRRRRRRRRRRRRRRRRRkRJH_C0M,NMRRRRRR--TCkH0NRhhBR5R_wuh2qh
RRRRRRRRRRRRRRRRRRRRRRRRCRMoM_HVR,RRRRRRR--hNCo0CHPRVHMH0MH$BR5R_wuQQhwh Qa2R
RRRRRRRRRRRRRRRRRRRRRRMRRCMo_FNslDR,RR-R-RoMCNP0HCFRMsDlNH8xCRMMFxFCs
RRRRRRRRRRRRRRRRRRRRRRRRCRMoC_8MlFsNRD,RR--MNCo0CHPRM8CFNslDCHx8wR5uz_1A)hmv2qp
RRRRRRRRRRRRRRRRRRRRRRRRCRMoC_xsRF,RRRRRR---5jRBuRw_)Z mR2
RRRRRRRRRRRRRRRRRRRRRRRRb_F#xFCs,RRRR-RR-jR+RR5BwZu_ 2)m
RRRRRRRRRRRRRRRRRRRRRRRRFRb#C_8MlFsNRD,RR--uHF#0CHPRM8CFNslDCHx8wR5uz_1A)hmv2qp
RRRRRRRRRRRRRRRRRRRRRRRRFRb#F_MsDlN,RRRRR--bHF#0CHPRsMFlHNDxRC8MxFMC
sFRRRRRRRRRRRRRRRRRRRRRRRRR#bF_VHM,RRRRRRR-b-RF0#HHRPCHHMVM$H0
RRRRRRRRRRRRRRRRRRRRRRRR#RHGR2;RRRRRRRRRR--ND0RC0N#RCFMRbHMkH0R#MRk	IMFMR

RR--a#EHRV8CCCss8FROMN#0MI0RHRDD0DCDRk$FRRHV0RECb	NONRoCL$F8RRH##0$MEHC#xDNLCR
R-F-RslRHblDCCCM08#RNRNsCDkRMlsLC#R3
RMOF#M0N0bRVE#8D$EM0__FssDCNRA:Rm mpqRh;RR--8CCVs8sCRMOF#M0N0R

RR--)kC0sRM#0RECO#DN#ERIHROEXNRVDRD#HFM0
VRRk0MOHRFMB#DN#RVb5R
RRRRGRRRRRRRRRRR:z h)1emp V7_D0FN;RRRRRRRRRRRR-RR-DRVFHN0MboRF0HMRbHMkR0
RORRE	CO_sCsF:sRRmAmph qRR:=VNDF0E_OC_O	CFsssR2R-O-RE	CORsVFRsCsF
s#RRRRskC0sPMRN8DH_#Vb0CN0;R

RR--q0sHE0lCHVORk0MOH#FM,ER0CR#CFsbCNs0F#FR8R0MFRJsCkCHsRsbNN0lCC3s#
VRRk0MOHRFM"#NL"NR5s:oRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR-R"RRs5NoRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0
;
R-R-RCaE#NCRDIDF#ER0CNRL#lCRNR0EVOkM0MHF#FR0RCk#RC0ERV8CN0kDRDPNk
C#R-R-RRFV0HECsNRbsCNl0#Cs3aRRERk#0$ECRR8FVDkDR Q  DRVFHN0MboRF0HM3R

RMVkOF0HM+R""RRR5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HM-R""RRR5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HM*R""RRR5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HM/R""RRR5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMsR"CRl"5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMlR"FR8"5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0
;
R-R-R#ANHbORNlsNCs0CR#DH0R
R-s-RF8kM_$#0D-CRRD1CC#O0RC0ERksFMM8HoDRNoHFs0REl0kFR#RC
RR--oskN8RR-CsG0NHRL0N#R888CRR0F0RECCRM8H0VREFCRbNCs0MHFRR0FNR88bOsCHF#HMR
R-O-RE	CO_sCsF-sRRCWEMVR"NCD#"kR0sRM#FRVVhRqhNRM8FsPCVIDFRCOEO
	#R-R-RM8CFNslDCHxRW-RERCM"DVN#RC"0Mks#VRFVCR8MlFsNMDRkClLssRbF#OC#oHM
R
RVOkM0MHFR8N8RR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0kRoNRs8RRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#;RR--MLklCFsRVkRoNRs8L#H0
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFM#0kLs0NORR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0kRoNRs8RRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#;RR--MLklCFsRVkRoNRs8L#H0
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFMl0kDH$bDRR5
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0kRoNRs8RRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#;RR--MLklCFsRVkRoNRs8L#H0
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFM8HHP85CR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0oskN8RRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H0;-RR-kRMlsLCRRFVoskN8HRL0R#
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN;R

RMVkOF0HMCRslMNH8RCs5R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0
;
RkRVMHO0FlMRFD8kF
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0Mo0Rk8NsRRRRR:RRRahqzp)qRRRR:V=RD0FN_NoksL8_H;0#R-R-RlMkLRCsFoVRk8NsR0LH#R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF;N0
R
R-s-RCbOHsNFODR
RVOkM0MHFROsCHFbsORND5R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0
;
RkRVMHO0F8MRH8PHCbL$.
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0Mo0Rk8NsRRRRR:RRRahqzp)qRRRR:V=RD0FN_NoksL8_H;0#R-R-RlMkLRCsFoVRk8NsR0LH#R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF;N0
R
R-v-RkHD0bRD$NkOOlNkD0RCRskC#D=0RRsD*RO+R
VRRk0MOHRFMlRNO5R
RR,RDRRs,ORRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0
;
R-R-Rk1JNRsCs0FFRD5ND6R(cNRL#RC8HDlbCMlC0HN0FRM#M8CCRH0E#R2
RMVkOF0HMJR#s50R
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRRRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0D
C;RRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFMQh#_C0oNHRPC5oNsRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm ;qh
R
R-----------------------------------------------------------------------------R
R-O-RFNlbsVCRk0MOH#FM
-RR-,R=R,/=R,>=R,<=RR<,>l,RNlGHkRl,lHHMl
kl
VRRk0MOHRFMC5JRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-JRCkRND=R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpq:hR=DRVF_N0OOEC	s_Cs;Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm Rqh:V=RD0FN_M8CFNslDCHx2R
RRCRs0MksRmAmph q;R

RMVkOF0HMCRMRR5RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--MRF0CNJkD=R/
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpq:hR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMApmm ;qh
R
RVOkM0MHFRRD05RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-D-RCR##0MENRR<
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm Rqh:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMmRAmqp h
;
RkRVMHO0FoMR0RR5RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCosNs0CRN0EM
R>RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp h=R:RFVDN80_CsMFlHNDx
C2RRRRskC0sAMRm mpq
h;
VRRk0MOHRFMD5CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-CRD#0#RERNMFCsRJDkNRR0F<R=
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm Rqh:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMmRAmqp h
;
RkRVMHO0FoMRCRR5RRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RCosNs0CRN0EMsRFRkCJN0DRF=R>
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpq:hR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMApmm ;qh
R
R-h-RCRC80FFRPDCsFRN80REC8NCVkRD0P#CsH#FMRRFV0#ECCR
RVOkM0MHFR""=RDR5,RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0F"MR/R="5RD,sRR:z h)1emp V7_D0FN2CRs0MksRmAmph q;R
RVOkM0MHFR=">"DR5,RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0F"MR<R="5RD,sRR:z h)1emp V7_D0FN2CRs0MksRmAmph q;R
RVOkM0MHFR"">RDR5,RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0F"MR<R"R5RD,sRR:z h)1emp V7_D0FN2CRs0MksRmAmph q;R

RMVkOF0HM?R"=R"R5RD,sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5,RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R">R"R5RD,sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5,RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtBR;
RMVkOF0HM?R"<R"R5RD,sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5,RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB
;
RkRVMHO0F#MR0l8_NE0OR,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp hR;
RMVkOF0HMHRVMs8_H0oEl0F#Rs5NoRR:z h)1emp V7_D0FN;RR$:aR17p_zmBtQ2R
RRCRs0MksRaQh )t ;R
RVOkM0MHFRMVH8C_DVF0l#50RNRso:hRz)m 1p7e _FVDNR0;$RR:1_a7ztpmQ
B2RRRRskC0sQMRhta  
);RkRVMHO0FlMRNlGHk5lRDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRMlHHllkR,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;
-RR-FROMsPC#MHFRMVkOF0HMR#
RR--BPFMC#s0RCFMRFVDNM0HoFRbHRM0MLklCHsRMR0FN0MFE3Cs
R
RVOkM0MHFR#sCHRxC5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRwFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRCOEOC	_sssFRRRR:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNH_xCH:MRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx;-RR-#RzC RQ C RGM0C8RC8wRu
RORRF0M#NRM08FCMsDlNHRxCR:RRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFMsHC#x5CR
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFwDNM0HoFRbHRM0HkMb0R
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0EROC_O	CFsssRRRRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHx_RHM:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR;R-z-R#QCR R  CCG0M88CR
wuRRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF;N0
R
RVOkM0MHFR_0FVNDF0Rd.5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;R
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0EROC_O	CFsssRRRRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHx_RHM:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR;R-z-R#QCR R  CCG0M88CR
wuRRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VFdN0.
;
RkRVMHO0F0MRFD_VFnN0c
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRRRR:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFsR:RRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDxHC_MRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0;nc
R
RVOkM0MHFR_0FVNDF0U4.RR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;
RORRF0M#NRM0sMFk80_#$RDCR:RRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsFRsRRRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;Fs
RRRRMOF#M0N0CR8MlFsNxDHCM_HRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC;RR--zR#CQ   R0CGCCM88uRw
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN4;.U
R
R-B-RFCMPsR0#NVMRbMRH0NFRMpR1eMR5CCC88FRVs$R#MC0E#2H#
VRRk0MOHRFM0#F_D5PRNRso:hRz)m 1p7e _FVDNR02skC0s1MRap7_mBtQ_Be a;m)
NRRD#HNR_0F1p08FOoHe0COFHsR#FR0_P#DRhrz)m 1p7e _FVDNs0RCs0kMaR17m_pt_QBea Bm;)9
NRRD#HNR_0F1_08pHFoOC_eOs0FRRH#0#F_DrPRz h)1emp V7_D0FNR0sCkRsM1_a7pQmtB _eB)am9
;
R-R-RMBFP0Cs#MRNRRVbHFM0RRNM#_08koDFHPO_CFO0s#R5k2DP
VRRk0MOHRFM0#F_kRDP5oNsRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQeB_ mBa)R;
RHNDN0#RF0_18FzpoeHOCFO0s#RHR_0F#PkDRhrz)m 1p7e _FVDNs0RCs0kMaR17p_zmBtQ_Be a9m);R
RNNDH#FR0_810_Fzpo_HOe0COFHsR#FR0_D#kPzRrh1) m pe7D_VFRN0skC0s1MRaz7_pQmtB _eB)am9
;
R-R-R8#0_FkDo_HOP0COF0sRFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:1_a7ztpmQeB_ mBa)R;
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=VNDF0G_CbCFMMI0_HE80;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RsRRCs0kMhRz)m 1p7e _FVDN
0;
-RR-MRQ0CCosFR0RFVDNR0
RMVkOF0HMFR0_FVDN50R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRQ:Rhta  
);RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)pRRRRR:=VNDF0G_CbCFMMI0_HE80;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRRRR:V=RD0FN_NVsOF0HMH_I8;0ER-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$2DCR-R-RksFMM8HobRF0MHF
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--sDCNRR0FVNDF0R
RVOkM0MHFR_0FVNDF0
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR: R)q
p;RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)pRRRRR:=VNDF0G_CbCFMMI0_HE80;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRRRR:V=RD0FN_NVsOF0HMH_I8;0ER-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--kHM#o8MCRR0FVNDF0R
RVOkM0MHFR_0FVNDF0
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7R;
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC2RR--sMFk8oHMR0FbH
FMRRRRskC0szMRh1) m pe7D_VF;N0
R
R-#-RHCoM8FR0RFVDNR0
RMVkOF0HMFR0_FVDN50R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)RqpR:RR=DRVF_N0CFGbM0CM_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azqRpRR=R:RFVDNV0_s0NOH_FMI0H8ER;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRksFM#8_0C$DRRRR:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR2R-s-RF8kMHRMoFHb0FRM
RsRRCs0kMhRz)m 1p7e _FVDN
0;
-RR-MRk#MHoCV8RH8GCRHbFM00RFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-k-RMo#HMRC8VCHG8FRbHRM0HkMb0R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)RqpR:RR=DRVF_N0CFGbM0CM_8IH0RE;RR--I0H8EVRFRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--I0H8EVRFRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCk#RCHCCGRC0#CMH#FM
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--#MHoCV8RH8GCRHbFM00RFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHM
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--sMFk8oHMR0FbH
FMRRRRskC0szMRh1) m pe7D_VF;N0
R
R-#-RH_xCsRC#VOkM0MHF#R
R-Q-RMo0CC0sRFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRRaQh )t ;R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR2R-s-RF8kMHRMoFHb0FRM
RsRRCs0kMhRz)m 1p7e _FVDN
0;
-RR-CRsN0DRFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRRq) pR;
R#RRH_xCsRC#RRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--kHM#o8MCRR0FVNDF0R
RVOkM0MHFR_0FVNDF0
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7h_z1hQt 
7;RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$2DCR-R-RksFMM8HobRF0MHF
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--#MHoC08RFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 71hQt 
7;RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$2DCR-R-RksFMM8HobRF0MHF
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--#PkDRR0FVNDF0R
RVOkM0MHFR_0FVNDF0
R5RRRRNRsoRRRRR1:Raz7_pQmtB _eB)am;R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2
RsRRCs0kMhRz)m 1p7e _FVDN
0;
-RR-MRk#MHoCV8RH8GCRHbFM00RFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;RR--kHM#o8MCRGVHCb8RF0HMRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHM
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCk#RCHCCGRC0#CMH#FM
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--#MHoCV8RH8GCRHbFM00RFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHC
8;RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-FRskHM8MFoRbF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0
;
R-R-RFVDN00RFMRk#MHoCR8
RMVkOF0HMFR0_#kMHCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRR:RRRahqzp)q;RRRR-R-RMDCoR0EFFVRkk0b0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF2-RR-EROCRO	VRFsCFsssR#
RsRRCs0kMhRz)m 1p7e _1zhQ th7
;
R-R-RFVDN00RFHR#o8MC
VRRk0MOHRFM0#F_HCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRR:RRRahqzp)q;RRRR-R-RMDCoR0EFFVRkk0b0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF2-RR-EROCRO	VRFsCFsssR#
RsRRCs0kMhRz)m 1p7e _t1Qh; 7
R
R-b-RkFsb#RC:BPFMC#s0RVNRD0FNRR0FkHM#o8MCRGVHCb8RF0HM
VRRk0MOHRFM0kF_VCHG8
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VHbRM0bk
RRRRMOF#M0N0CRDVH0_MG8CRRRRRQ:Rhta  R);RR--HCM0oRCsb0Ns
RRRRMOF#M0N0HRso_E0HCM8GRRRRQ:Rhta  R);RR--VOsN0MHFRsbN0R
RRFROMN#0MF0RPVCsD_FI#D0$CRR:VCHG8P_FCDsVF#I_0C$D_b0$C=R:RGVHCF8_PVCsD_FI#D0$CR;R-#-RNs0kN
0CRRRRO#FM00NMRksFM#8_0C$DRRRR:HRVG_C8sMFk80_#$_DC0C$bRRRR:V=RH8GC_ksFM#8_0C$D;-RR-FRskHM8MRo
RORRF0M#NRM0OOEC	s_CsRFsR:RRRmAmph qRRRRRRRRRRRRRRRRR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhRRRRRRRRRRRRRRRRR=R:RFVDN80_CsMFlHNDx
C2RRRRskC0szMRh1) m pe7V_kH8GC;R

RR--VNDF0FR0Ro#HMRC8VCHG8FRbH
M0RkRVMHO0F0MRFV_#H8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RbMRHb
k0RRRRO#FM00NMRVDC0M_H8RCGRRRR:hRQa  t)R;R-H-RMo0CCbsRN
s0RRRRO#FM00NMRosHEH0_MG8CRRRR:hRQa  t)R;R-V-Rs0NOHRFMb0Ns
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;-RR-NR#0Nks0RC
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0MO0RE	CO_sCsFRsRRRR:Apmm RqhRRRRRRRRRRRRRRRRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRRRRRRRRRRRRRRRRRRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMhRz)m 1p7e _H#VG;C8
R
R-#-RH_xCsRC#P#CsH#FM
-RR-DRVFRN00kFRMo#HM
C8RkRVMHO0F0MRFM_k#MHoC58R
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7R;
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR2R-O-RE	CORsVFRsCsF
s#RRRRskC0szMRh1) m pe7h_z1hQt 
7;
-RR-DRVFRN00#FRHCoM8R
RVOkM0MHFR_0F#MHoC58R
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRR:hRz)m 1p7e _t1Qh; 7
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs2FsR-R-RCOEOV	RFCsRsssF#R
RRCRs0MksR)zh p1me_ 71hQt 
7;
-RR-kRbs#bFCB:RFCMPsR0#NDRVFRN00kFRMo#HMRC8VCHG8FRbH
M0RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RbMRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8
RRRRMOF#M0N0PRFCDsVF#I_0C$DRV:RH8GC_CFPsFVDI0_#$_DC0C$bRR:=VCHG8P_FCDsVF#I_0C$D;-RR-NR#0Nks0RC
RORRF0M#NRM0sMFk80_#$RDCR:RRRGVHCs8_F8kM_$#0D0C_$RbCR:RR=HRVG_C8sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0MO0RE	CO_sCsFRsRRRR:Apmm RqhRRRRRRRRRRRRRRRRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRRRRRRRRRRRRRRRRRRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMhRz)m 1p7e _HkVG;C8
R
R-V-RD0FNRR0F#MHoCV8RH8GCRHbFMR0
RMVkOF0HMFR0_H#VGRC85R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-bRVRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7#GVHC
8;RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DCR-R-R0#Nk0sNCR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0DRC;RR--sMFk8oHM
RRRRMOF#M0N0EROC_O	CFsssRRRRA:Rm mpqRhRRRRRRRRRRRRRRRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRRRRRRRRRRRRRRRR:V=RD0FN_M8CFNslDCHx2R
RRCRs0MksR)zh p1me_ 7#GVHC
8;
-RR-DRVFRN00sFRC
NDRkRVMHO0F0MRFC_sN5DR
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsM)p q;R

RR--VNDF0FR0R0HMCsoC
VRRk0MOHRFM0HF_Mo0CC5sR
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR2R-O-RE	CORsVFRsCsF
s#RRRRskC0sQMRhta  
);
-RR-FRwsCResFHDoFROl0bNNDLHH
0$RkRVMHO0FsMRC0NDF0LH#NR5s:oRRq) ps2RCs0kMaR17p_zmBtQ_Be a;m)
VRRk0MOHRFML#H00CFsN5DRNRso:aR17p_zmBtQ_Be a2m)R0sCkRsM)p q;R

RR--v#NbR0lCNoDFHDONRDPNk
C#RkRVMHO0F0MRF4_jRR5
RNRRsRoR:hRz)m 1p7e _FVDNR0;RRRRRRRRR-RR-DRVFHN0MboRF0HMRbHMkR0
RXRRvRqu:aR17m_ptRQB:'=Rj
'2RRRRskC0szMRh1) m pe7D_VF;N0
R
RVOkM0MHFR_Q#XNR5sRoRRRR:z h)1emp V7_D0FN2CRs0MksRmAmph q;R
RVOkM0MHFR_0FXRj45oNsRRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMFR0_4XjZNR5s:oRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F0MRFX_zj54RNRso:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VF;N0
R
R-a-RECC#RF0IRFbsOkC8sRC#ICCsRbOFHRC8FRk0F0VRELCRFR8$LNCOkR#C0$ECRFbsP
C8R-R-RsPC$#RkCDVkRsVFRMPC8RFs#ObCHOVHRoNDF0sHE8lRCDPCFCblMR0
RR--ANsC	k_MlsLCRMOFP0Cs#RRNVNDF0oHMRHbFMM0RkClLsMRH0HFR0R'#b0Ns#R
R- -RGMbFCRM0HL#RHCN#8$RLR
-4
bRRsCFO8CksRCLsNM	_kClLs
R5RRRRNRsoRRRRRRRR:MRHRhRz)m 1p7e _FVDN
0;RRRR8FCMsDlNHRxC:MRHRmRAmqp h=R:RFVDN80_CsMFlHNDx
C;RRRROOEC	s_CsRFs:MRHRmRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRVOsN0RRRRRRR:kRF0hRz)m 1p7e _1zhQ th7R;
RCRRGMbFRRRRR:RRR0FkR)zh p1me_ 71hQt R7;RR--h ma:qRR848RRR0FoRC00RECsDCNRbCGFMMC0R!
R#RRHRoMRRRRR:RRR0FkR71a_mzpt2QB;R

RFbsOkC8sLCRs	CN_lMkLRCs5R
RRsRNoRRRRRRRRRR:HRMRz h)1emp V7_D0FN;R
RRCR8MlFsNxDHCRR:HRMRApmm Rqh:V=RD0FN_M8CFNslDCHx;R
RREROC_O	CFsssRR:HRMRApmm Rqh:V=RD0FN_COEOC	_sssF;R
RRsRVNRO0RRRRRRR:FRk0z h)1emp k7_VCHG8R;R-N-RRlMkLRCsLIC0CRCM4R3jNRM8.
3jRRRRCFGbMRRRRRRR:kRF0hRz)m 1p7e _t1Qh; 7R-R-Rahm R:RqR884FR0R0oCRC0ERNsCDGRCbCFMM
0!RRRR#MHoRRRRRRRR:kRF0aR17p_zmBtQ2
;
R-R-RshFlHNDx0CRN#	CRVNRs0NOHRFMNRM8NRM8CFGbM0CMR8NMRMOFP0Cs#ER0CHlRM
0FR-R-RVNRD0FNHRMobMFH0kRMlsLC37RRFRC#0REC#VEH0oHMR8NMRC0ERksFMM8HoR3
RR-- FGbM0CMRRH#Nk##lRC80LFRCHRLN8#CRRL$-
4
RkRVMHO0FMMRFNslDCHxRR5
RVRRs0NORRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;-RR-sRVNHO0FRM,kFMMsDlNH8xC
RRRRbCGFRMRRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;RRR-C-RGMbFCRM0-,R4RsMFlHNDx
C8RRRR#MHoRRRRRRRRRRRRRRRRRRRR:aR17p_zmBtQ;RRRRRRRR-R-Ro#HMHRL0R
RR0R#H$O	RRRRRRRRRRRRRRRRRRR:1_a7ztpmQ:BR=jR''R;R-1-R0	HO$HRL0sR5F8kMH2Mo
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azqRpRR=R:RFVDNC0_GMbFC_M0I0H8ER;R-#-RHRxCFFVRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRRRR:V=RD0FN_NVsOF0HMH_I8;0ER-R-Rx#HCVRFR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR;R-z-R#QCR R  CCG0M88CR
wuRRRRO#FM00NMRkMoNRs8RRRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H02RRR-o-Rk8NsR0LH#R
RRCRs0MksR)zh p1me_ 7VNDF0
;
R-R-Rb GFMMC0#RHR#N#k8lCRR0FLLCRHCN#8$RLR
-4RkRVMHO0FMMRFNslDCHxRR5
RVRRs0NORRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;R-R-R#kMHCoM8HRVGRC8bMFH0R
RRGRCbRFMRRRRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;RRR--CFGbM0CMR4-R,FRMsDlNH8xC
RRRRo#HMRRRRRRRRRRRRRRRRRRRR1:Raz7_pQmtBR;RRRRRR-RR-HR#oLMRHR0
R#RR0	HO$RRRRRRRRRRRRRRRR:RRR71a_mzptRQB:'=RjR';RR--1O0H	L$RH50RsMFk8oHM2R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)RqpR:RR=DRVF_N0CFGbM0CM_8IH0RE;RR--#CHxRRFVFbk0kC0RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)pRRRRR:=VNDF0s_VNHO0FIM_HE80;-RR-HR#xFCRVkRF00bkRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC;RR--zR#CQ   R0CGCCM88uRw
RRRRMOF#M0N0oRMk8NsRRRRRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R2RRR--oskN8HRL0R#
RsRRCs0kMhRz)m 1p7e _FVDN
0;
VRRk0MOHRFMMlFsNxDHC
R5RRRRVOsN0RRRRRRRRRRRRRRRRz:Rh1) m pe7h_z1hQt R7;R-RR-MRk#MHoCR8
RCRRGMbFRRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh; 7RRRRR-R-RbCGFMMC0RR-4M,RFNslDCHx8R
RRHR#oRMRRRRRRRRRRRRRR:RRR71a_mzpt;QBR-R-Ro#HMHRL0R
RR0R#H$O	RRRRRRRRRRRRR:RRR71a_mzptRQB:'=RjR';RR--1O0H	L$RH50RsMFk8oHM2R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRR--k8#CRsVFRx#HHRMoF$MD
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0MM0RoskN8RRRR:RRRahqzp)qRRRR:V=RD0FN_NoksL8_H20#R-RR-kRoNRs8L#H0
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR-- FGbM0CMRRH#Nk##lRC80LFRCHRLN8#CRRL$-R4
RMVkOF0HMFRMsDlNHRxC5R
RRsRVNRO0RRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHCR8;RRRRRR--kHM#o8MCRGVHCb8RF0HM
RRRRbCGFRMRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;RRRRR-C-RGMbFCRM0-,R4RsMFlHNDx
C8RRRR#MHoRRRRRRRRRRRRRRRRR1:Raz7_pQmtBR;R-#-RHRoML
H0RRRR#O0H	R$RRRRRRRRRRRRRR1:Raz7_pQmtB=R:R''j;-RR-0R1H$O	R0LHRF5skHM8M
o2RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-RR-#RkCV8RF#sRHMxHoMRFDR$
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR;R-z-R#QCR R  CCG0M88CR
wuRRRRO#FM00NMRkMoNRs8RRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R2RRR--oskN8HRL0R#
RsRRCs0kMhRz)m 1p7e _FVDN
0;
-RR-PRFCFsDN88CRsPC#MHF#R
RVOkM0MHFR""+R5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR+R"RRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""+R5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR+R"RRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""-R5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR-R"RRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""-R5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR-R"RRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""*R5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR*R"RRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""*R5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR*R"RRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""/R5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR/R"RRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFR""/R5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MR/R"RRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRC"sl5"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRs"ClRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRC"sl5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRs"ClRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRF"l85"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRl"F8RR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRF"l85"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRl"F8RR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R

RR--FsPCD8FNCO8RFNlbsVCRk0MOH#FM
VRRk0MOHRFM"R="RDR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksRmAmph q;R
RVOkM0MHFR="/"5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMmRAmqp hR;
RMVkOF0HM>R"=R"R5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpRRRRskC0sAMRm mpq
h;RkRVMHO0F"MR<R="RR5D:hRz)m 1p7e _FVDNR0;sRR:)p q2RRRR0sCkRsMApmm ;qh
VRRk0MOHRFM"R>"RDR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksRmAmph q;R
RVOkM0MHFR""<R5RRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMmRAmqp hR;
RMVkOF0HM=R""RRR5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0RRRRskC0sAMRm mpq
h;RkRVMHO0F"MR/R="RR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMApmm ;qh
VRRk0MOHRFM"">=RDR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksRmAmph q;R
RVOkM0MHFR="<"5RRDRR:)p q;RRs:hRz)m 1p7e _FVDNR02RsRRCs0kMmRAmqp hR;
RMVkOF0HM>R""RRR5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0RRRRskC0sAMRm mpq
h;RkRVMHO0F"MR<R"RRR5D: R)qRp;sRR:z h)1emp V7_D0FN2RRRR0sCkRsMApmm ;qh
VRRk0MOHRFM"R="RDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksRmAmph q;R
RVOkM0MHFR="/"5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMmRAmqp hR;
RMVkOF0HM>R"=R"R5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  R)2skC0sAMRm mpq
h;RkRVMHO0F"MR<R="RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsMApmm ;qh
VRRk0MOHRFM"R>"RDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksRmAmph q;R
RVOkM0MHFR""<R5RRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMmRAmqp hR;
RMVkOF0HM=R""RRR5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0F"MR/R="RR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm ;qh
VRRk0MOHRFM"">=RDR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksRmAmph q;R
RVOkM0MHFR="<"5RRDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp hR;
RMVkOF0HM>R""RRR5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0F"MR<R"RRR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm ;qh
VRRk0MOHRFM""?=RDR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) pR2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?=RDR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2RRCRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?=RDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?=RDR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?/"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?>RDR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?>"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM""?<RDR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
VRRk0MOHRFM"=?<"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzpt;QB
-RR-HRlMkHllMRN8NRlGkHllPRFCFsDN
8#RkRVMHO0FlMRNlGHk5lRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRHlMHk5lRDRR:z h)1emp V7_D0FN;RRs: R)qRp2RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRNlGHk5lRDRR:)p q;RRs:hRz)m 1p7e _FVDNR02RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRHlMHk5lRDRR:)p q;RRs:hRz)m 1p7e _FVDNR02RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRNlGHk5lRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRHlMHk5lRDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRNlGHk5lRDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FlMRHlMHk5lRDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;----------------------------------------------------------------------------
-RR-FRDoNHODkRVMHO0F
M#R-R--------------------------------------------------------------------------
-
RkRVMHO0F"MRM"F0RDR5RRRR:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFM"8NM"5RRDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRs"F"RRR5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMMR"N"M8R,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRM"FsRDR5,RRs:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFM"sGF"5RRDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRM"GFRs"5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0R;
RR--e0COFNsRM#8R0k8_DHFoOkRVMHO0F,M#Rl#NC#RNRMVkOF0HMH#RMkRMlHCsO0_#8R
RVOkM0MHFRM"N85"RDRR:1_a7ztpmQRB;sRR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMNR"MR8"5:DRR)zh p1me_ 7VNDF0s;RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRFRs"5:DRR71a_mzpt;QBR:sRR)zh p1me_ 7VNDF0R2
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRFRs"5:DRR)zh p1me_ 7VNDF0s;RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRM8NM"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7D_VF2N0
RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRN"MMR8"5:DRR)zh p1me_ 7VNDF0s;RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRM"FsRR5D:aR17p_zmBtQ;RRs:hRz)m 1p7e _FVDN
02RRRRskC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFM"sMF"DR5Rz:Rh1) m pe7D_VF;N0R:sRR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRF"Gs5"RDRR:1_a7ztpmQRB;sRR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMGR"FRs"5:DRR)zh p1me_ 7VNDF0s;RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0F"MRGsMF"DR5R1:Raz7_pQmtBs;RRz:Rh1) m pe7D_VF2N0
RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRM"GFRs"5:DRR)zh p1me_ 7VNDF0s;RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDN
0;R-R-R8)CkHO0FFMRbNCs0#Fs,NR#lNCR#kRMlHCsO0_#8kRVMHO0F
M#RkRVMHO0F"MRN"M8RDR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRM8NM"DR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRFRs"RDR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRM"FsRDR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRG"FsRDR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;RkRVMHO0F"MRGsMF"DR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQ
B;
-RR-FRh0RC:"N#D"",R#"sN,#R"D,D"RD"#sR","DsF"MRN8sR"FRs"MRF0HDlbCMlC03C8
R
R-----------------------------------------------------------------------------R
R-)-RClOFl8CMCw8Rk0MOH#FMRFVslER0C RQ ( R6qcRbMbC8
HGR-R--------------------------------------------------------------------------
--
-RR-CRs0Mks#RRGIEH0RC0ERo#HMVRFR
$3RkRVMHO0FBMRF#b$HRoM5RG,$RR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0
;
R-R-R0)Ck#sMR*$RR*.*MFRVsMRH0sCoNPDRNCDk#VRFRIhRHF0EkO0RFklb0oHMR*.*MR
RVOkM0MHFRN1OD5LR
RRRRR$RRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RhRRRRRRRRRRRRRRRRRRRRRR:hRQa  t)R;RR-RR-GRCbCFMM00RF8RN8RRRRR
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF;N0
R
R-)-RCs0kM$#RR.*R*R*MVRFsHCM0oDsNRDPNkRC#FhVRR0IHE0FkRlOFbHk0M.oR*
*MRkRVMHO0F1MROLNDRR5
R$RRRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRRhRRRRRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;RRRRR-C-RGMbFCRM00NFR8R8RRRR
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN;R

RR--skC0sRM#0RECkHMLN8#CRbCGFMMC0VRFRRG
RMVkOF0HMFRpo5LRGRR:z h)1emp V7_D0FN2CRs0MksRaQh )t ;R
RVOkM0MHFRopFLGR5Rz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp 17_Q th7
;
R-R-R0sCk#sMRC0ERGMC0CRsb#sCCNM0LRDCMoCHEsLFRRFVGMRHRC0ERs8HCHO0F0MRFsIN8
R$RkRVMHO0FhMRCNG0Vs0CRR5
RGRR,RR$RRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm Rqh:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp h=R:RFVDN80_CsMFlHNDx
C2RRRRskC0szMRh1) m pe7D_VF;N0
R
R-)-RCs0kMa#R)Rz HXVRRRH#ksMF8CCs8HRI0YER3R
RVOkM0MHFRFzMss8CC58RG$,RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm ;qh
VRRk0MOHRFMwHHM05CRGRRRRRRR:hRz)m 1p7e _FVDNR02skC0sAMRm mpq
h;RkRVMHO0FQMR#MMNRR5GRRRRR:RRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h
;
R-R-RMwkOF0HMFR0R0sCkRsMO#FM00NM#R3
RMVkOF0HMCRxsbFVRR5
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=VNDF0G_CbCFMMI0_HE80;-RR-GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802-RR-sRVNHO0FRM
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FMMRNbMVRR5
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=VNDF0G_CbCFMMI0_HE80;-RR-GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802-RR-sRVNHO0FRM
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FJMRMVNMb
R5RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;R-C-RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RFVDNV0_s0NOH_FMI0H8ER2R-V-Rs0NOH
FMRRRRskC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFMb_F#HVMVb
R5RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;R-C-RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RFVDNV0_s0NOH_FMI0H8ER2R-V-Rs0NOH
FMRRRRskC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFMM_CoHVMVb
R5RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;R-C-RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RFVDNV0_s0NOH_FMI0H8ER2R-V-Rs0NOH
FMRRRRskC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFMM_CoxFCsV5bR
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq:pR=DRVF_N0CFGbM0CM_8IH0RE;RR--CFGbM0CM
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=DRVF_N0VOsN0MHF_8IH0RE2RR--VOsN0MHF
RRRR0sCkRsMz h)1emp V7_D0FN;R
R-#-RH_xCsRC#P#CsH#FM
VRRk0MOHRFMxFCsV5bR
RRRRx#HCC_s#RR:z h)1emp V7_D0FN2RRRRRRRRR--PHNsNCLDRRH#F$MDRCk#RsVFRx#HH
MoRRRRskC0szMRh1) m pe7D_VF;N0
VRRk0MOHRFMMVNMb
R5RRRR#CHx_#sCRz:Rh1) m pe7D_VF2N0RRRRRRRR-P-RNNsHLRDCHF#RMRD$kR#CVRFs#HHxMRo
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FJMRMVNMb
R5RRRR#CHx_#sCRz:Rh1) m pe7D_VF2N0RRRRRRRR-P-RNNsHLRDCHF#RMRD$kR#CVRFs#HHxMRo
RsRRCs0kMhRz)m 1p7e _FVDN
0;RkRVMHO0FbMRFH#_MbVVRR5
R#RRH_xCsRC#:hRz)m 1p7e _FVDNR02RRRRR-RR-NRPsLHNDHCR#MRFDk$R#VCRF#sRHMxHoR
RRCRs0MksR)zh p1me_ 7VNDF0R;
RMVkOF0HMCRMoM_HVRVb5R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RsPNHDNLC#RHRDFM$#RkCFRVsHR#xoHM
RRRR0sCkRsMz h)1emp V7_D0FN;R
RVOkM0MHFRoMC_sxCFRVb5R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RsPNHDNLC#RHRDFM$#RkCFRVsHR#xoHM
RRRR0sCkRsMz h)1emp V7_D0FN;-

-NbsoRlN#0$MEHC##V_FV-
-RDs0_M#$0#ECHF#RV
V
R-R-=========================================================================
==R-R-Rs#0HRMoNRM800CGHwFRk0MOH#FM
-RR-===========================================================================
R
R-I-RsCH0#:R1    :wwwwwwwwR
RbOsFCs8kC)RWQRa 5R
RRRRpRRRRRRRR:MRHFRk0p Qh;RRRRRRRRRRRR-RR-ORNO#C#Rb0$CbR5F0HMC
s2RRRRezqp RRRRRR:HRMRRhRz)m 1p7e _FVDNR0;RR--PkNDCFR0RHIs0RC
RKRRzQ1aw7Q RH:RMRRRR71Q :RR=HRso;E0RRRR-I-REEHOR8#HCFR0R#[k0$HVRG0C0R
RRQRw Rp7RRRR:MRHRRRRWaQ7]=R:R;j2RRRRR-RR-HRI8R0EFVVRH8CD
R
R-)-RC#N8R 1  w wwwwwwRw,"R3"NRM8"R:"NRsCHFoMs
C8RsRbF8OCkRsC)7 qRR5pR:RRRFHMkp0RQ;h Rpeqz: RR0FkR)zh p1me_ 7VNDF0
2;RsRbF8OCkRsC)7 qRR5pR:RRRFHMkp0RQ;h Rpeqz: RR0FkR)zh p1me_ 7VNDF0R;
RRRRRRRRRRRRRRRRRmtm7RR:FRk0RmRAmqp h
2;
NRRD#HNR A)qH7R# R)qr7Rp Qh,hRz)m 1p7e _FVDNR0,Apmm 9qh;R
RNNDH#)RA Rq7H)#R Rq7rhpQ z,Rh1) m pe7D_VF9N0;R
RNNDH#WRA) QaRRH#Wa)Q pRrQ,h R)zh p1me_ 7VNDF01,RQ,7 R7WQa;]9
NRRD#HNRhAQq_)Y)7 qRRH#)7 qRQrphR ,z h)1emp w7_pamq,mRAmqp h
9;RDRNHRN#AqQh))Y_ Rq7H)#R Rq7rhpQ z,Rh1) m pe7p_wm9qa;R
RNNDH#QRAhYq)_QW)aH R#)RWQRa rhpQ z,Rh1) m pe7D_VF,N0R71Q W,RQ]7a9
;
RsRbF8OCkRsCmQW)a5 R
RRRRRpRRRRRR:RRRFHMkp0RQ;h RRRRRRRRRRRRR-R-RONOCR##0C$bRF5bHCM0sR2
ReRRq pzRRRRRH:RMRRRR)zh p1me_ 7VNDF0R;R-P-RNCDkRR0FI0sHCR
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHER0;R-RR-ERIHROE#CH8RR0F[0k#HRV$00CG
RRRR wQpR7RR:RRRRHMRWRRQ]7aRR:=jR2;RRRRR-R-R8IH0FERVHRVC
D8
-RR-ORm0RNDs8CNR0IHENRb8M8HoM,RFCR#bNNs0#FsRCk#8R
RbOsFCs8kC)Rm Rq75RpRRRR:HkMF0QRphR ;ezqp RR:FRk0z h)1emp V7_D0FN2R;
RFbsOkC8smCR)7 qRR5pR:RRRFHMkp0RQ;h Rpeqz: RR0FkR)zh p1me_ 7VNDF0R;
RRRRRRRRRRRRRRRRRmRtm:7RR0FkRARRm mpq;h2
NRRD#HNRamBq)p_ Rq7Hm#R)7 qRQrphR ,z h)1emp w7_pamq,mRAmqp h
9;RDRNHRN#mqBap _)qH7R#)Rm Rq7rhpQ z,Rh1) m pe7p_wm9qa;R
RNNDH#BRma_qpWa)Q #RHR)mWQRa rhpQ z,Rh1) m pe7p_wm,qaR71Q W,RQ]7a9
;
R-R-RG]CRHIs0ICRHR0Eb8N8H,MoRRMF#NCbsFN0sR#
RFbsOkC8s]CRWa)Q 
R5RRRRpRRRRRRRRRR:HkMF0QRphR ;RRRRRRRRRRRRRR--NCOO#0#R$RbC5HbFMs0C2R
RRqRepRz RRRR:MRHRRRRz h)1emp V7_D0FN;-RR-NRPDRkC0IFRsCH0
RRRR1KzaQQw :7RRRHMR1RRQR7 RR:=sEHo0R;RR-R-RHIEO#ERHR8C0[FRkH#0V0$RC
G0RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2R;RRRRRRR--I0H8EVRFRCVHD
8
R-R-RG]CRNsC8HRI0bERNH88MRo,M#FRCsbNNs0F##RkCR8
RFbsOkC8s]CR)7 qRR5p:MRHFRk0p Qh;qRepRz :kRF0hRz)m 1p7e _FVDN;02
bRRsCFO8CksR ])q57RpRRRRH:RM0FkRhpQ e;Rq pzRF:Rkz0Rh1) m pe7D_VF;N0
RRRRRRRRRRRRRRRRRRRt7mmRF:RkR0RRmAmph q2R;
RHNDN]#R )X_ Rq7H]#R)7 qRQrphR ,z h)1emp w7_pamq,mRAmqp h
9;RDRNHRN#]_ X)7 qRRH#]q) 7pRrQ,h R)zh p1me_ 7wqpma
9;RDRNHRN#]_ XWa)Q #RHR)]WQRa rhpQ z,Rh1) m pe7p_wm,qaR71Q W,RQ]7a9
;
R-R-RDs0_M#$0#ECHF#RMR
R-s-bNNolRM#$0#ECHF#_MR
R
-RR-CRs0Mks#1R":    w:wwwwww
w"RkRVMHO0F0MRF0_#soHMRN5PDRkC:hRz)m 1p7e _FVDNR02skC0s1MRah)QtR;
RHNDNa#Rm1_Aah)Qt#RHR_am1Qa)hrtRz h)1emp w7_pamqR0sCkRsM1Qa)h;t9
NRRD#HNR_amAqQh)1Y_ah)Qt#RHR_am1Qa)hrtRz h)1emp w7_pamqR0sCkRsM1Qa)h;t9
R
R-)-RCs0kMN#RRX] Rs#0H,MoR0IHENRb8M8HoR
RVOkM0MHFR_0FEs#0HRMo5DPNk:CRR)zh p1me_ 7VNDF0s2RCs0kMaR1)tQh;R
RNNDH#mRa_X] _)1aQRhtHa#Rm1_]ah)QtzRrh1) m pe7p_wmRqaskC0s1MRah)Qt
9;
-RR-CR)0Mks#MRN8ORF0RND#H0sMRo,IEH0R8bN8oHM
VRRk0MOHRFM0FF_#H0sM5oRPkNDCRR:z h)1emp V7_D0FN2CRs0MksR)1aQ;ht
NRRD#HNR_ammqBapa_1)tQhRRH#amm_1Qa)hrtRz h)1emp w7_pamqR0sCkRsM1Qa)h;t9
R
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoRRRRRRRRRRRRRR:RRR)1aQ;htR-RR-HRLM$NsRs#0H
MoRRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802R
RRCRs0MksR)zh p1me_ 7VNDF0R;
RHNDNV#Rs_FlLs#0HRMoHV#Rs_Fl#H0sMroR1Qa)hRt,hzqa),qpRahqzp)q
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7VNDF0
9;RDRNHRN#VlsF_MLHN_s$#H0sMHoR#sRVF#l_0MsHo1Rrah)Qth,Rq)azqRp,hzqa)
qpRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _FVDN;09
VRRk0MOHRFMVlsF_0F#soHMRR5
RFRR#H0sMRoRRRRRRRRRRRRRR:RRR)1aQ;htR-RR-ORm0RND#H0sMRo
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=VNDF0G_CbCFMMI0_HE80;R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820E
RRRR0sCkRsMz h)1emp V7_D0FN;R
RNNDH#sRVFFl_OD0N_s#0HRMoHV#Rs_FlFs#0HRMor)1aQ,htRahqzp)q,qRhaqz)pR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp V7_D0FN9
;
RkRVMHO0FVMRs_FlEs#0HRMo5R
RR#RE0MsHoRRRRRRRRRRRRRRRRRR:1Qa)hRt;R-R-RGECRs#0H
MoRRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802R
RRCRs0MksR)zh p1me_ 7VNDF0R;
RHNDNV#Rs_FlE_CG#H0sMHoR#sRVFEl_#H0sMroR1Qa)hRt,hzqa),qpRahqzp)q
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRs0MksR)zh p1me_ 7VNDF0
9;
VRRk0MOHRFMVlsF_s#0HRMo5R
RR#RL0MsHo:RRR)1aQ;htRRRRRRRRRRRRRRRRR-R-RMLHNRs$#H0sMRo
R#RRH_xCsRC#:hRz)m 1p7e _FVDNR02RRRRR-RR-#RkCV8RF#sRHMxHoMRFD
$RRRRRskC0szMRh1) m pe7D_VF;N0
NRRD#HNRFVsl#_L0MsHo#RHRFVsl0_#soHMRar1)tQh,hRz)m 1p7e _FVDNR0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRskC0szMRh1) m pe7D_VF9N0;R
RNNDH#sRVFLl_HsMN$0_#soHMRRH#VlsF_s#0HRMor)1aQ,htR)zh p1me_ 7VNDF0R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0sCkRsMz h)1emp V7_D0FN9
;
RkRVMHO0FVMRs_FlFs#0HRMo5R
RR#RF0MsHo:RRR)1aQ;htRRRRRRRRRRRRRRRRR-R-R0mON#DR0MsHoR
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RCk#8FRVsHR#xoHMRDFM$RR
RsRRCs0kMhRz)m 1p7e _FVDN
0;RDRNHRN#VlsF_0FON#D_0MsHo#RHRFVsl#_F0MsHo1Rrah)Qtz,Rh1) m pe7D_VF
N0RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _FVDN;09
R
RVOkM0MHFRFVsl#_E0MsHo
R5RRRREs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-E-RC#GR0MsHoR
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RCk#8FRVsHR#xoHMRDFM$RR
RsRRCs0kMhRz)m 1p7e _FVDN
0;RDRNHRN#VlsF_GEC_s#0HRMoHV#Rs_FlEs#0HRMor)1aQ,htR)zh p1me_ 7VNDF0R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRCs0kMhRz)m 1p7e _FVDN;09
M
C8NRbOo	NCDRVF_N0oCCMs_HOb;	o
N
bOo	NCFRL8V$RD0FN_MoCCOsH_ob	R
H#
-RR-kRq0sEFRP7NHA8RHF#Eb8R5LEH#F@b@PDE83oFs2R
R-----------------------------------------------------------------------------R
R-0-R$RbC8DCON0sNH#FM
-RR----------------------------------------------------------------------------
R
R-a-RERH#8CCVs8sCRMOF#M0N0HRID0DRCRDD$RFkH0VREbCRNNO	oLCRFR8$H##R$EM0Cx#HNCLD
-RR-sRFRbHlDCClM80CRRN#sDCNRlMkL#Cs,CR#0FR0Rs"0kRC"H#VR$EM0Cx#HNCLD3R
RO#FM00NMREVb8$D#M_0EFss_CRND:mRAmqp h=R:Rk0sCR;R-8-RCsVCsRC8O#FM00NM
R
R-0-R$#bCRRFVLMFk8$NsRMOF8HH0F
M#R$R0bLCRF8kMN_s$0C$bRRH#5sMFl,NDRVHMH0MH$x,RC,sFRM8CFNslD
2;
-RR-kRMDsDRNCMoRsNsNO$RF0M#N
M0RFROMN#0Mh0RqRwu:hRz)m 1p7e _FVDN50RjFR8IFM0RR42RR:=5EF0CRs#='>Rj;'2
ORRF0M#NRM0he1pR1:Raz7_pQmtB _eB)amRR5j8MFI04FR2=R:R05FE#CsRR=>'2j';R

RR--1ObCHRNDP#CsHRFMF"VRlHHMl"klRR0F8#FRFRlCLMFk8$NsRCOEOM	HoR
RVOkM0MHFRMlHCpR5,RR):hRQa  t)R2
RsRRCs0kMhRQa  t)#RH
LRRCMoHR-R-RMVkOF0HMHRlMkHllR
RRVRHRR5p=hRQa  t)F'DIsRFR=)RRaQh )t 'IDF2ER0CRM
RRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRR&RR"zFMLkCM88kRMlsLCR#bN#,C8R#INRDNRHs0CNkDR#?C8"R
RRRRRRCR#PHCs0C$RsssF;R
RRRRRskC0sjMR;R
RRMRC8VRH;R
RRCRs0MksRMlHHllkR,5pR;)2
CRRMV8Rk0MOHRFMlCHM;R

RR--tCCMsCN0#ER0CNRL#MCRkClLsFRVsER0CGRCbCFMMM0RFNslDNHx0MHFRVFV#3C0
VRRk0MOHRFMo_CMCFGbMN_L#5CR
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq
p2RRRRskC0s1MRQ th7R
RHR#
RPRRNNsHLRDCskC#D:0RRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2
LRRCMoH
RRRR#sCkRD0RRRRRRRRRRRRRRRRR:RR=FR50sEC#>R=R''42R;
RsRRCD#k0CR5GMbFC_M0I0H8E2-4RR:=';j'
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0FoMRCCM_GMbF_#LNC
;
R-R-R0QMCsoCRsPC#MHFRRFV0REC"oDF.O"RFNllM58RO0FMskHL0RC8Lu$RCs0CREq#CCM8MR2
RMVkOF0HMFRDo5.RqRR:hzqa)2qpR0sCkRsMhzqa)RqpHR#
RPRRNNsHLRDCJ0kFH0CMRh:Rq)azq
p;RRRRPHNsNCLDR#sCkRD0RRR:hzqa)Rqp:j=R;R
RLHCoMR
RRkRJFC0HM:0R=RRq/;R.
RRRRHIEDJCRkHF0CRM0>RRjDbFF
RRRRJRRkHF0CRM0:J=RkHF0CRM0/;R.
RRRRsRRCD#k0RRR:s=RCD#k0RR+4R;
RCRRMD8RF;Fb
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0FDMRF;o.
R
R-w-Rk0MOHRFM#HHlDRNs00FREQCRpAmtRMVkOF0HMMRHRavq] _)qRp
RMVkOF0HMFRDo5.RqRR:)p q2CRs0MksRaQh )t R
H#RRRRPHNsNCLDR:YRRq) pR;
RPRRNNsHLRDChRR:Q hatR ):j=R;R
RLHCoMR
RRVRHRR5q=3R4jsRFR=qRRjj32ER0CRM
RRRRR0sCkRsMjR;
RCRRMH8RVR;
RYRRRR:=qR;
RHRRVR5q>3R4j02RE
CMRRRRRERIHRDCY=R>Rj.3RFDFbR
RRRRRRRRY:Y=RR./R3
j;RRRRRRRRh=R:R+hRR
4;RRRRRMRC8FRDF
b;RRRRRCRs0MksR
h;RRRRCRM8H
V;RRRR-m-RRY<RR4<R
RRRRHIEDYCRR4<R3DjRF
FbRRRRRRRY:Y=RR.*R3
j;RRRRRRRh:h=RR4-R;R
RRMRC8FRDF
b;RRRRskC0shMR;R
RCRM8VOkM0MHFRoDF.
;
R-R-RsbkbCF#:CRa#00RELCRF8kMNRs$O8FMHF0HMF#RVRRN)DCNRlMkL
CsRsRbF8OCkRsC00C#_kLFMs8N$
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:MRHRq) pR;RR-RR-MRQb,k0RMOFP0CsC08RFCRsNRD
RORRF0M#NRM0VOsN0MHF_8IH0:ERRRHMhzqa);qpR-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERR:HhMRq)azqRp;RR--DoCM0FERVuRwRbCGFMMC0R
RRFROMN#0M80RCsMFlHNDxRCRRRR:HAMRm mpq:hR=sR0kRC;RR--zR#CQ   R0CGCCM88uRw
RRRRsPNHDNLC0RL$RbC:kRF0FRLkNM8s0$_$;bC
RRRRsPNHDNLCFRDoR.H:kRF0hRQa  t)R
RRRR2HR#
RORRF0M#NRM0CFGbMN_L#:CRRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0RRj2:R=
RRRRRMoC_bCGFLM_N5#CCFGbM0CM_8IH0;E2R-RR-GRCbCFMMF0RVCV#0R
RRFROMN#0MC0RGlb_H:MRRt1QhR 75R4.8MFI0jFR2=R:
RRRR-RR5#sCH5xCCFGbMN_L#RC,42d2R4+R;RRRRR--vHHMlRklMlFsNCDRGMbFC
M0RRRRO#FM00NMRbCG_0CG_MlHR1:RQ th74R5.FR8IFM0RRj2:R=
RRRRRbCG_MlHRV-Rs0NOH_FMI0H8ER;RRRRRR-RR-HRvMkHllFRVsCR8MlFsNCDRGMbFC
M0RRRRPHNsNCLDRoDF.oNsRQ:Rhta  R);RRRRRRRR-D-RFRo.FNVRslokC
M0RCRLoRHMRR--VOkM0MHFR#0C0F_LkNM8sR$
R-RR-ERBCRO	0#FRCHCRVER0CGRCbCFMMH0R#HRLoMRCFEko
RRRRR--hCF0RN0E0ER0CsRNoCklMH0R#DRNI#N$RRNMNFL#DCk0RDPNkNCR0ER0Hb#RF0HM3R
RRFRDos.No=R:RoDF.s5No
2;RRRRHNVRs=oRRjj3RC0EMR
RRRRRLb0$C=R:RsxCFR;
RCRRDV#HRbCGFMMC0H_I8R0E>4R4RC0EMRRRR-RR-GR bCFMMV0RF)sRCRNDH4#R4nR5cHRL0R2
RRRRR$L0b:CR=FRMsDlN;R
RRDRC#RC
RRRRRRHVD.FoNRso<FR0_0HMCsoC5bCG_MlH2ER0CRM
RRRRRHRRVCR8MlFsNxDHCER0CRM
RRRRRRRRRRHVD.FoNRso<FR0_0HMCsoC5bCG_0CG_MlH2ER0CRM
RRRRRRRRRLRR0C$bRR:=xFCs;R
RRRRRRRRRCCD#
RRRRRRRRRRRR$L0b:CR=CR8MlFsN
D;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRRRHVD.FoNRso<FR0_0HMCsoC5bCG_MlH2R-40MEC
RRRRRRRRRRRR$L0b:CR=CRxs
F;RRRRRRRRRDRC#RC
RRRRRRRRRLRR0C$bRR:=MlFsNRD;RRRRRRRRRRRRRR--BRNM#D0HDCRsb#sCCRM00#EHRlMkL
CsRRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R
RRRRRCHD#VGRCbCFMMI0_HE80R4<R4ER0CRM
RRRRRHRRVFRDos.NoRR>0HF_Mo0CCCs5GMbF_#LNC42+RC0EMR
RRRRRRRRRLb0$C=R:RVHMH0MH$R;
RRRRRCRRD
#CRRRRRRRRR0RL$RbC:M=RFNslDR;
RRRRRCRRMH8RVR;
RRRRR#CDCR
RRRRRR0RL$RbC:M=RFNslDR;
RRRRR8CMR;HV
RRRR8CMR;HV
RRRRoDF.:HR=FRDos.NoR;
R8CMRFbsOkC8s0CRC_#0LMFk8$Ns;R

RR--bbksF:#CRk)FMR8#8CCbMM8HoMRFRC0ERN#00FCRVER0CsR"F8kM_$#0D
C"R-R-RopFH0ORNM	CRFVslR
R-"-RW0ENRC PsB$RFklb0RCs1COHM#0H0ER1F8kDRFiMILRqFRk0wNDF0oHMRHuFMq0RsEH0lHC0OR"
RR--L7$RN8PHRDtF8sLCo4R5g2g4
VRRk0MOHRFMOOEC	F_skRM85R
RRsRVN_O0HRMRRRRRRRRRR:RRR71a_mzpt;QBR-R-RbHMkV0Rs0NOH
FMRRRR#MHoRRRRRRRRRRRRRRRRR1:Raz7_pQmtBR;R-#-RHRoML
H0RRRRsNClHCM8sRRRRRRRRRRRRz:Rht1Qh; 7RRRR-s-RCHlNMs8CRR0FsMFk8sRVFRl
R#RR0	HO$RRRRRRRRRRRRRRR:aR17p_zmBtQRR:=';j'RRRRR-R-RH10OR	$L
H0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$CR2R-s-RF8kMHRMo0C$b
RRRR0sCkRsMApmm 
qhR#RH
RRRRsPNHDNLCCRs#0kDRRRRRA:Rm mpq
h;RRRRPHNsNCLDR_FsskC8ORC8:aR17p_zmBtQ;R
RLHCoM-RR-kRVMHO0FOMRE	CO_ksFMR8
RsRRCD#k0=R:RDVN#
C;RRRRH5VRsNClHCM8sC'DMEo0Rj>R2ER0CRMRRRRR-H-RVCRslMNH8RCsHNMRRDMkDsRNs
N$RRRRRsRF_8sCk8OCRR:=F5sRsNClHCM8sRR&#O0H	;$2
RRRRsRRF8kMH_MoOCN#RO:RNR#CsMFk80_#$RDCHR#
RRRRRIRRERCMsMFk8C_MN#sC0>R=RRRRRRRRR-RR-FR)kRM8hsCNC,#0RV8CN0kDR8lFCR
RRRRRRRRRHsVRCHlNMs8C5lsCN8HMCEs'H2oER'=R40'RERCMRR--sMFk8R
RRRRRRRRRRVRHRC5slMNH8'CsDoCM0>ERRR420MEC
RRRRRRRRRRRRHRRV5R5F5sRsNClHCM8sC5slMNH8'CsEEHo-R4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0sFRCHlNMs8C'IDF2=2RR''4
RRRRRRRRRRRRRRRRRRRF#sR0	HO$RR='24'
RRRRRRRRRRRRRRRRFRRssRVN_O0H=MRR''42ER0CRM
RRRRRRRRRRRRR-RR-NRv	0CRELCRFF00lHRL0CRxsHFRVFRb#L#HDHCRVCRIRCNsRRN04
/.RRRRRRRRRRRRRRRRskC#D:0R=sR0k
C;RRRRRRRRRRRRRMRC8VRH;R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRR#sCkRD0:5=RVOsN0M_HR'=R4F'Rs0R#H$O	R'=R4;'2
RRRRRRRRRRRR8CMR;HV
RRRRRRRRCRRMH8RVR;
RRRRRIRRERCMsMFk8M_HV>R=RRRRRRRRRRRRR-RR-FRskRM8kHbRVFRb#HH0PRC,CCD#Rk0sM0ONCR3
RRRRRRRRRRHVFss_CO8kC=8RR''4R8NMRo#HMRR='Rj'0MEC
RRRRRRRRRRRR#sCkRD0:0=Rs;kC
RRRRRRRRCRRMH8RVR;
RRRRRIRRERCMsMFk8C_MoVHMRR=>RRRRR-RR-FRskRM88MFIRRHVMNCo0CHP,DRC#0CRsOkMN30C
RRRRRRRRHRRVsRF_8sCk8OCR'=R4N'RM#8RHRoM=4R''ER0CRM
RRRRRRRRRsRRCD#k0=R:Rk0sCR;
RRRRRRRRR8CMR;HV
RRRRRRRRCIEMFRsk_M8xFCsRR=>RRRRRRRRRRRRRR--sMFk8FR0I8NsRRjRRkasM0ONCR
RRRRRRRRRMDkD;R
RRRRRCRM8OCN#RksFMM8HoN_O#
C;RRRRCRM8H
V;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMEROC_O	sMFk8
;
R-R-RsbkbCF#:FR)k#M8Rb8CCHM8MFoRMER0C0R#NR0CF0VRE"CRsMFk80_#$"DC
-RR-MRk#MHoCP8RCHs#FRM
RFbsOkC8sVCRbF_skRM85R
RRsRVN_O0HRMR:MRHRhRz1hQt R7;RRRRRRRRR-R-RbHMkV0Rs0NOH
FMRRRRCFGbMM_HRRR:HRMR1hQt R7;RRRRRRRRRRRR-H-RM0bkRbCGFMMC0R
RRsRVN_O0FRk0:kRF0hRz1hQt R7;RRRRRRRRR-R-R0FkbRk0VOsN0MHF
RRRRbCGFFM_k:0RR0FkRt1Qh2 7RRH#RRRRRRRRRR--Fbk0kC0RGMbFC
M0RCRLoRHMRR--bOsFCs8kCbRV_ksFMR8
RHRRVMRN8VR5s0NO_2HMR'=R40'RERCMRRRRR-RR-sRwNHO0FHMR#DRND4R""R
RRRRRCFGbMk_F0=R:RbCGFHM_MRR+4R;
RRRRRNVsOF0_k:0R=FR0_#kMHCoM8,5jRNVsOF0_kE0'H+oE4
2;RRRRCCD#
RRRRCRRGMbF_0FkRR:=CFGbMM_H;R
RRRRRVOsN0k_F0=R:RNVsOH0_MRR+4R;
RCRRMH8RVR;
R8CMRFbsOkC8sVCRbF_sk;M8
R
R-a-RERH#P#CsHRFMFLVRs	CN_lMkLRCs8#FCMR'0ODNDRD"ONV##bR"
RFbsOkC8sLCRs	CN_lMkLRCs5RRRRRRRRRRRR-RR-MRH0MCsNPDRCHs#FRM
RNRRsRoRRRRRR:RRRRHMR)zh p1me_ 7VNDF0R;
RVRRbb0$RRRRR:RRRRHMRDPNHV8_bN#00
C;RRRR8FCMsDlNHRxC:MRHRmRAmqp h=R:Rk0sCR;
RVRRs0NORRRRR:RRR0FkR1zhQ th7R;
RCRRGMbFRRRRR:RRR0FkRt1Qh2 7R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:Rs-NoF'DIR;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RoNs'oEHER;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRO#FM00NMRbCGFLM_NR#CRRRR:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2RjR
:=RRRRRCRoMG_Cb_FMLCN#5bCGFMMC0H_I820E;RRR-C-RGMbFCRM0F#VVCR0
RPRRNNsHLRDCCRGb:QR1t7h RG5Cb'FMsoNMC
2;RCRLo
HMRRRRVOsN0VR5s0NOH_FMI0H8ER-48MFI0jFR2=R:
RRRRzRRht1QhR 75_0F#5DPN5so-84RF0IMFVR-s0NOH_FMI0H8E222;R
RRsRLCON	NR#C:NRO#VCRbb0$R
H#RRRRRERICbMRFx#_CRsF|CRMoC_xs=FR>R
RRRRRRsRVNRO05NVsOF0HMH_I820ERR:=';j'
RRRRRRRRbCGRRRRRRRRRRRRRRRRRRRR:-=RCFGbMN_L#
C;RRRRRERICbMRF8#_CsMFlRND|CRMoC_8MlFsN=DR>R
RRRRRRVRHRM8CFNslDCHxRC0EMR
RRRRRRRRRCRGbRRRRRRRRRRRRRRRRR:RR=CR-GMbF_#LNCR;
RRRRRRRRRNVsO50RVOsN0MHF_8IH0RE2:'=Rj
';RRRRRRRRCCD#
RRRRRRRRCRRGRbRRRRRRRRRRRRRRRRRR=R:RG-Cb_FMLCN#R4-R;R
RRRRRRRRRVOsN0VR5s0NOH_FMI0H8E:2R=4R''R;
RRRRRCRRMH8RVR;
RRRRRCIEMFRb#F_MsDlNRM|RCMo_FNslDRR|b_F#HRMV|CRMoM_HV>R=
RRRRRRRRNVsO50RVOsN0MHF_8IH0RE2:'=R4
';RRRRRRRRCRGbRRRRRRRRRRRRRRRRR:RR=QR1t7h 5oNs5bCGFMMC0H_I8-0E4FR8IFM0R2j2;R
RRRRRRGRCbCR5GMbFC_M0I0H8E2-4RR:=MRF0C5GbCFGbM0CM_8IH04E-2R;
RRRRRCIEM0RFE#CsR
=>RRRRRRRRNC##sh0Rmq_W)hhQtR
RRRRRRRRRsFCbsw0Rpamq_ht  B)Q_tui'#HM0ONMCN_MlRC
RRRRRRRRR"&RAq) iz_hv)A :RR"&R
RRRRRRRRR"0vCN0R#NR0C8CC0O80CRRHMVLb_s	CN_lMkLRCsbOsFC"##
RRRRRRRR#RRCsPCHR0$IMNsH;Mo
RRRRRRRRR--ObFlDCC0RC0ER#ONCH,RVRRNhRqho#FCR,HMRhNRqOhRF#lCR0Fk3R
RRRRRRGRCbRRRRRRRRRRRRRRRRRRRRR:=5EF0CRs#='>R4;'2
RRRRRRRRNVsO50RVOsN0MHF_8IH0RE2:'=R4
';RRRRCRM8OCN#RCLsNN	O#
C;RRRRCFGbM=R:RbCG;R
RCRM8bOsFCs8kCsRLC_N	MLklC
s;
-RR-kRbs#bFCV:RD0FNHRMobMFH0FR0R1zhQ th7R
R-z-R#RC8L0$RFM_H0CCos0,RFM_k#MHoCR8,NRM80#F_HCoM8kRVMHO0F
M#RsRbF8OCkRsCVNDF0F_0_#kMHCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRH:RMzRRh1) m pe7D_VF;N0RRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRPHNsNCLDRo#HMRRRRRRRRF:Rk10Raz7_pQmtBR;RRRRRRRRR-#-RHRoMFFVRkk0b0R
RRNRPsLHNDVCRsRNORRRRR:RRR0FkR1zhQ th7R;RRRRRRRRRR-R-R#kMHCoM8HRLN8#CR0Fkb
k0RRRRO#FM00NMRM8CFNslDCHxRH:RMARRm mpqRh;RRRRRRRRRRRR-0-RkRsMF8MRCsMFlHNDxHN0FRM
RORRF0M#NRM0L#HNRRRRRRRR:MRHRqRhaqz)pR;RRRRRRRRRR-RR-HRLNV#RFVsRH8GCRHbFMR0
RORRF0M#NRM0sMFk80_#$RDC:MRHRFRsk_M80C$b2#RHRRRRR-RR-FRskHM8MloRCF0E8R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:Q hatR ):-=RlCHM5oNs'IDF,sRNoF'DIR2;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0GRCbCFMMI0_HE80RQ:Rhta  :)R=sRNoH'EoRE;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRsPNHDNLCsRVNRO0RRRRRRRRRz:Rht1QhR 75NVsON'sM2oC;-RR-MRH0MCsNPDRCHs#FFMRVsRVNRO
RPRRNNsHLRDCHo#HMRRRRRRRR:RRR71a_mzpt;QBRRRRRRRRR-RR-MRH0MCsNPDRCHs#FFMRVHR#oRM
RPRRNNsHLRDCCRGbRRRRRRRRR:RRRaQh )t ;-RR-GR bCFMMR0
RPRRNNsHLRDCCFGbMRRRRRRRR:RRRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2R-R-ROeC0HFsxRC8C
GbRRRR-A-RNR#C08FRH8PHCsRVNHO0FLMR$R
RRNRPsLHNDVCRs_NO#VEH0RRRRRR:zQh1t7h Rs5VNEO'H+oEdFR8IFM0R;j2R-R-RNwsOF0HMER#HCV08R
RRNRPsLHND#CRE0HVRRRRRRRRRRR:Q hat; )
RRRRsPNHDNLCCRslMNH8RCsRRRRRz:Rht1QhR 758.RF0IMF2Rj;R
RRNRPsLHNDsCRF8kMRRRRRRRRRRR:1_a7ztpmQRB;RRRRRRRRR-R-RksFMA8RQRa
RoLCHRM
RHRR#MHoRRRRRRRRRRRRRRRRR:RR=FR0_4Gj5oNs5oNs'oEHE;22
RRRRR--CFGbM0CMRR/=',j'RsMFlRNDVNDF0oHMRHbFMR0
RCRRGMbFRRRRRRRRRRRRRRRRR:RR=FR0_5j41hQt N75s5oRCFGbM0CM_8IH04E-RI8FMR0Fj,22R''X2R;
RCRRGMbF5bCGFMMC0H_I8-0E4:2R=FRM0GRCb5FMCFGbM0CM_8IH04E-2R;
RCRRGRbRRRRRRRRRRRRRRRRRR:RR=FR0_0HMCsoCRG5Cb2FM;R
RR-R-RowHkRsCFRk00RECVOsN0MHF
RRRRNVsOR0RRRRRRRRRRRRRRRRRRR:=5EF0CRs#='>Rj;'2RRRRRR--VDHDR0IHECRxsRF
RVRRs0NORs5VN'O0EEHo2RRRR:RR=4R''R;RR-RR-8Rq8ER0C4R"33j"
RRRRH#EVR0RRRRRRRRRRRRRRRRRRR:=5NVsOE0'H-oE4-2RRbCG;R
RRVRHRNVsOF0HMH_I8R0E>sRVN'O0EEHoRC0EMRRRRRRRRRRRR-R-RMBNRDFM$#RkCHR#x.C-R0LH#R
RRRRRVOsN0VR5s0NO'oEHER-48MFI0jFR2=R:R1zhQ th70R5FD_#PNR5s-o54FR8IFM0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVR-s0NO'oEHE222;R
RRDRC#RCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-RMONRCk#RDNDR0LH#R
RRRRRVOsN0VR5s0NO'oEHER-48MFI0VFRs0NO'oEHEs-VNHO0FIM_HE802=R:
RRRRRRRR1zhQ th70R5FD_#PNR5s-o54FR8IFM0Rs-VNHO0FIM_HE802;22
RRRR8CMR;HV
RRRRNVsOE_#HRV0:V=Rs0NOR"&Rj"jj;R
RRVRHRH#EV<0RR0jRERCMRRRRRRRRRRRRRRRRR-R-RCmPsFVDIR
RRRRRVOsN0=R:R05FE#CsRR=>'24';R
RRDRC#RC
RRRRRNVsOE_#HRV0:#=RE0HV_osHE50RVOsN_H#EVR0,#VEH0
2;RRRRRsRVNRO0RRRRRR:=VOsN_H#EV50RVOsN_H#EVE0'HRoE8MFI0dFR2R;
RRRRRlsCN8HMCRsR:V=Rs_NO#VEH0.R5RI8FMR0Fj
2;RRRRR-R-RksFM58RsMFk8C_xsIFRHRDDLN$b#0#RERH#NRM80MskOCN02R
RRRRROCN#RksFM#8_0C$DR
H#RRRRRRRRIMECRksFMM8_CCNs#=0R>R
RRRRRRRRRsMFk8=R:RlsCN8HMC.s52MRN8R
RRRRRRRRRRRRRRRRRRs5VNRO05Rj2F5sRF5sRsNClHCM8s4R5RI8FMR0Fj2222R;
RRRRRIRRERCMsMFk8M_HV>R=
RRRRRRRRsRRF8kMRR:=sNClHCM8s25.R8NMR0MFRHH#o
M;RRRRRRRRIMECRksFMM8_CMoHV>R=
RRRRRRRRsRRF8kMRR:=sNClHCM8s25.R8NMRHH#o
M;RRRRRRRRIMECREF0CRs#=R>
RRRRRRRRRksFM:8R=jR''R;
RRRRR8CMR#ONCR;
RRRRRRHVsMFk8RR='R4'0MEC
RRRRRRRRNVsO:0R=sRVNRO0+;R4
RRRRCRRMH8RVR;
RCRRMH8RVR;
RVRRsRNO:V=Rs0NO;R
RRHR#o:MR=#RHH;oM
CRRMb8RsCFO8CksRFVDN00_FM_k#MHoC
8;
-RR-kRbs#bFCs:RCs0kMN#RRsbN0VRFRPNRCFO0s0,RERH#VOkM0MHFRRH#ECCsROLCNCk#
-RR-sRFRs5VNsO0RF50_0HMCsoC5H#EV20GRI8FMR0Fj;22
-RR-NROMR'0L#CR$EM0Cx#HCH8RMFR#l#CR$EM0C##HRF0FD
#3RkRVMHO0F#MRlDNDVOsN0
R5RRRRNRsoRRR:zQh1t7h ;R
RRER#HRV0:qRhaqz)pR2
RsRRCs0kMaR17p_zmBtQ
HRR#R
RRNRPsLHNDFCRs:GRR71a_mzpt;QB
LRRCMoH
RRRRGFsRR:=N5so#VEH0
2;RRRRVRFsHMRHRoNs'MsNoDCRF
FbRRRRRVRHR<HRRH#EV00RE
CMRRRRRRRRFRsG:N=RsHo52sRFRGFs;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RRCRs0MksRGFs;R
RCRM8VOkM0MHFRN#lDsDVN;O0
-RR-------------------------------------------------------------------------R-
RR--eHH#LRDCVOkM0MHF#R
R-------------------------------------------------------------------------
--
-RR-kRbs#bFCO:RFCMPsR0#0RECMNCo0CHPR8HMC0GRFRRNbHF#0CHPRCFM
-RR-CRMoHN0PHCRMO8HCN#RsHCRDoDCNHDRM4R4nNcRM48Rj3(ndR
RVOkM0MHFR_0F#PkDRR5
RNRRs:oRR)zh p1me_ 7VNDF0R2RRRRRRRRRR-RR-bRVROPC0
FsRRRRskC0s1MRaz7_pQmtB _eB)am
HRR#R
RRNRPsLHNDsCRCD#k0RR:1_a7ztpmQeB_ mBa)NR5sDo'C0MoER-48MFI0jFR2R;
RoLCHRMR-V-Rk0MOHRFM0#F_0k8_DHFoOC_POs0F
RRRRRHVN'soDoCM0<ERR04RE
CMRRRRRCRs0MksRph1eR;
RCRRMH8RVR;
RsRRCD#k0=R:R71a_mzpt_QBea Bm5)RN2so;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0#F_k;DP
R
R-B-RFCMPsR0#NVMRbMRH0NFRMzR1pRe
RMVkOF0HMFR0_P#DRs5NoRR:z h)1emp V7_D0FN2CRs0MksR71a_tpmQeB_ mBa)#RH
LRRCMoH
RRRR0sCkRsM0#F_kRDP5oNs2R;
R8CMRMVkOF0HMFR0_P#D;R

RR--bbksF:#CRsMFlHNDxRC#NDRVFHN0MboRF0HMRlMkL
CsR-R-RHaE#CRPsF#HM#RN#Ckl#MRNRM"k#MHoCR8"HkMb0HRI0RE
RMVkOF0HMFRMsDlNHRxC5R
RRsRVNRO0RRRRRRRRRRRRRRRRRRR:z h)1emp z7_ht1Qh; 7R-RR-sRVNHO0FRM,kFMMsDlNH8xC
RRRRbCGFRMRRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;RRR-C-RGMbFC,M0RsMFlHNDxRC8L-$R4R
RRHR#oRMRRRRRRRRRRRRRRRRRRRR:1_a7ztpmQRB;RRRRRRRR-#-RHRoMA
QaRRRR#O0H	R$RRRRRRRRRRRRRRRRR:aR17p_zmBtQRR:=';j'R-R-RH10OR	$LRH05ksFMM8HoR2
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-Rx#HCVRFR0FkbRk0CFGbM0CM
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azqRpRR=R:RFVDNV0_s0NOH_FMI0H8ER;R-#-RHRxCFFVRkk0b0sRVNHO0FRM
RORRF0M#NRM0sMFk80_#$RDCR:RRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0MM0RoskN8RRRRRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#2RR--oskN8HRL0R#
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDRs#VNRO0RRRR:hRz1hQt 57RVOsN0H'Eo8ERF0IMF2Rj;-RR-ER#HCV08sRVNHO0FRM
RPRRNNsHLRDCsNVsOR0RR:RRR1zhQ th7VR5s0NOH_FMI0H8ER-48MFI0jFR2R;RRR--VOsN0MHF
RRRRsPNHDNLCGRCbRRRRRRRR1:RQ th7CR5GMbFC_M0I0H8ER+48MFI0jFR2R;R-C-RGMbFC
M0RRRRPHNsNCLDRGsCbRRRRRRR:QR1t7h RG5CbCFMMI0_HE80+84RF0IMF2Rj;-RR-CRs#0kDRbCGFMMC0R
RRNRPsLHNDsCRCFGbMRRRRRR:zQh1t7h RG5CbCFMMI0_HE80-84RF0IMF2Rj;RRR-C-RGMbFC
M0RRRRPHNsNCLDR#sCkRD0RRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8ER2;RR--skC#DR0
RPRRNNsHLRDC#VEH0RsRR:RRRaQh )t ;RRRR-RR-ER#HRV0NklFMR0
RPRRNNsHLRDC#O0H	R$GR:RRR71a_mzpt;QBR-RR-CRPsF#HMVRFRH#0O
	$RRRRO#FM00NMRbCGFLM_NR#C:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2RjR
:=RRRRRCRoMG_Cb_FMLCN#5bCGFMMC0H_I820E;RRR-C-RGMbFCRM0F#VVCR0
RPRRNNsHLRDCsMFk8x,RCssFCR#,HsMVC:#RRmAmph q;R
RLHCoM-RR-kRVMHO0FMMRFNslDCHx
RRRRsxCF#sCRR:=V#NDCR;
RHRRMCVs#:RR=NRVD;#C
RRRRksFMR8RRR:=V#NDCR;
R#RRE0HVs:RR=HRVMD8_ClV0FR#05_0FjV45s0NO2',R4R'2RRRR-w-RHRM80RECV#Hs04R""R
RRRRRRRRRRRRRRV-Rs0NOH_FMI0H8ERR-MNoksR8;RR--#0kLs0NORC0ERMDCoR0EIICRN
M0RRRRCRGb:s=RCx#HCCR5GMbF,GRCbC'DMEo02RR+#VEH0
s;RRRRH5VRF5sRVOsN0=2RR''j2ER0CRMRRR--ZFCs
RRRRxRRCssFC:#R=sR0k
C;RRRRCHD#V5R5CRGb<-=RsHC#xCC5GMbF_#LNCC,RGDb'C0MoE42-2MRN8CR8MlFsNxDHCR2
RRRRRRFs5G5CbRR<-#sCH5xCCFGbMN_L#RC,C'GbDoCM0-E24N2RMM8RF80RCsMFlHNDxRC20MEC
RRRRHRRVCR5G>bR=sR-Cx#HCG5Cb_FMLCN#,GRCbC'DMEo02s-VNHO0FIM_HE80-
42RRRRRRRRNRM88FCMsDlNHRxC0MEC
RRRRRRRRbCGRRRR:-=RsHC#xCC5GMbF_#LNCC,RGDb'C0MoE42-;R
RRRRRRER#HsV0RR:=-_0FHCM0oRCs5bCGF+MRRbCGFLM_N2#C;-RR-CRMIER#H
V0RRRRRDRC#RCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-s-RCs0kMCRxsRF
RRRRRxRRCssFC:#R=sR0k
C;RRRRRMRC8VRH;R
RRDRC#RHV5bCGRC>RGMbF_#LNC2-4RC0EMRRRR-R-RVHMH0MH$R
RRRRRHsMVC:#R=sR0k
C;RRRRCRM8H
V;RRRRHxVRCssFC0#RE
CMRRRRRCRs#0kDRR:=xFCsV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRR#CDHHVRMCVs#ER0CRM
RRRRR#sCkRD0:b=RFH#_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRDRC#RC
RRRRRs#VNRO0:V=Rs0NORD#sRH#EV;0sRRRRR-RR-ER#H
V0RRRRRVRHRH#EVR0s>RRj0MEC
R--RRRRR#RR0	HO$:GR=0R#H$O	RRFs5RFs5NVsO50R#VEH04s-RI8FMR0Fj222;R
RRRRRR0R#H$O	G=R:RH#0OR	$F#sRlDNDVOsN0VR5s0NO,ER#HsV0-;42
RRRRCRRD
#CRRRRRRRR#O0H	R$G:#=R0	HO$R;
RRRRR8CMR;HV
RRRRHRRVoRMk8NsRj>RRC0EMR
RRRRRRFRskRM8:O=RE	CO_ksFM58R
RRRRRRRRVRRs0NO_RHMR=RR>VR#s0NORo5Mk8Ns2R,
RRRRRRRRRo#HMRRRRRRRRR=>#MHo,R
RRRRRRRRRsNClHCM8sRRR=#>RVOsN0o5Mk8Ns-84RF0IMF2Rj,R
RRRRRRRRR#O0H	R$RRRRR=#>R0	HO$
G,RRRRRRRRRFRsk_M8#D0$C>R=RksFM#8_0C$D2R;
RRRRR8CMR;HV
RRRRHRRVFRskRM80MEC
RRRRRRRR_VbsMFk8s5VN_O0HRMR=#>RVOsN0VR5s0NOH_FMI0H8E+-4MNoks88RF0IMFoRMk8Ns2R,
RRRRRRRRRRRRRRRRCFGbMM_HR>R=RbCG5GsCbN'sM2oC,R
RRRRRRRRRRRRRRVRRs0NO_0FkRR=>sNVsO
0,RRRRRRRRRRRRRRRRRbCGFFM_k=0R>CRsG;b2
RRRRCRRD
#CRRRRRRRRsNVsO:0R=VR#s0NORs5VNHO0FIM_HE80-M4+oskN8FR8IFM0RkMoN2s8;R
RRRRRRCRsGRbRRR:=C5GbsbCG'MsNo;C2
RRRRCRRMH8RVR;
RRRRRR--skC#DR0
RRRRRGsCbRFM:z=Rht1QhR 75GsCbG5CbCFMMI0_HE80-84RF0IMF2Rj2R;
RRRRRGsCbRFM5bCGFMMC0H_I8-0E4R2RRRRRRRRR:M=RFs0RCFGbMG5CbCFMMI0_HE80-;42
RRRRsRRCD#k0sR5CFGbMN'sM2oCRRRRRRRRRRRRR=R:R)zh p1me_ 7VNDF0C5sGMbF2R;
RRRRR#sCkRD05R-48MFI0-FRVOsN0MHF_8IH0RE2:z=Rh1) m pe7D_VF5N0sNVsO;02
RRRR8CMR;HV
RRRR#sCkRD05bCGFMMC0H_I820ERR:=#MHo;RRRRR--#MHoRaAQ
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0FMMRFNslDCHx;R

RR--bbksF:#CRsMFlHNDxRC#NDRVFHN0MboRF0HMRlMkL
CsR-R-RHaE#CRPsF#HM#RN#Ckl#RRN"HkVG"C8RbHMkR0
RMVkOF0HMFRMsDlNHRxC5R
RRsRVNRO0RRRRRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-k-RMo#HMRC8VCHG8FRbH
M0RRRRCFGbMRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh; 7R-R-RbCGFMMC0M,RFNslDCHx8$RLR
-4RRRR#MHoRRRRRRRRRRRRRRRRRRRR:aR17p_zmBtQ;RRRRRRRR-R-Ro#HMHRL0R
RR0R#H$O	RRRRRRRRRRRRRRRRRRR:1_a7ztpmQ:BR=jR''R;R-1-R0	HO$HRL0sR5F8kMH2Mo
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azqRpRR=R:RFVDNC0_GMbFC_M0I0H8ER;R-#-RHRxCFFVRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRRRR:V=RD0FN_NVsOF0HMH_I8;0ER-R-Rx#HCVRFR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR;R-z-R#QCR R  CCG0M88CR
wuRRRRO#FM00NMRkMoNRs8RRRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H02RRR-o-Rk8NsR0LH#R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RPRRNNsHLRDCNksoM:#RR1zhQ th7VR5s0NO'oEHERR+VOsN0MHF_8IH0+ERRkMoN
s8RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2=R:R05FE#CsRR=>'2j';R
RLHCoM-RR-kRVMHO0FMMRFNslDCHx
RRRRoNskRM#5oNsk'M#EEHoRI8FMR0FlHNGlRkl5oNsk'M#EEHo-NVsOD0'C0MoE,+4R2j2R
:=RRRRRhRz1hQt 57R0#F_D5PRVOsN0;22
RRRR#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>NksoM
#,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=C>RGMbF,R
RRRRRRRRRRRRRRRRRRRRRR#RRHRoMRRRRRRRRR>R=Ro#HMR,
RRRRRRRRRRRRRRRRRRRRRRRR#O0H	R$RRRRRR=RR>0R#H$O	,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRkMoNRs8RRRRRRRR=M>RoskN8
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFRMsDlNH;xC
R
R-b-RkFsb#RC:MlFsNxDHCN#RRFVDNM0HoFRbHRM0MLklCRs
RR--a#EHRsPC#MHFR#N#k#lCR"NRkGVHCR8"HkMb0HRI0NERRH"#xsC_CR#"HkMb0R
RVOkM0MHFRsMFlHNDx5CR
RRRRNVsOR0RRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-k-RMo#HMRC8VCHG8FRbH
M0RRRRCFGbMRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;-RR-GRCbCFMMR0,MlFsNxDHCL8R$4R-
RRRRo#HMRRRRRRRRRRRRRRRRRR:1_a7ztpmQRB;RR--#MHoR0LH
RRRRH#0OR	$RRRRRRRRRRRRRRR:1_a7ztpmQ:BR=jR''R;R-1-R0	HO$HRL0sR5F8kMH2Mo
RRRRx#HCC_s#RRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRR-k-R#RC8VRFs#HHxMFoRM
D$RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC;RR--zR#CQ   R0CGCCM88uRw
RRRRMOF#M0N0oRMk8NsRRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#2R-R-RNoksL8RH
0#RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=#R-H_xCs'C#D;FI
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq:pR=HR#xsC_CE#'H;oE
RRRRsPNHDNLCCRs#0kDRRRRRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLCsRNo#kMRz:Rht1QhR 75NVsOE0'HRoE+sRVNHO0FIM_HE80RM+RoskN8R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RCRLoRHMRR--VOkM0MHFRsMFlHNDxRC
RNRRsMok#NR5sMok#H'Eo8ERF0IMFNRlGkHllNR5sMok#H'EoVE-s0NO'MDCo+0E4j,R2:2R=R
RRRRRzQh1t7h RF50_P#DRs5VN2O02R;
RsRRCD#k0=R:RsMFlHNDx5CRVOsN0RRRRRRRR=RR>sRNo#kM,R
RRRRRRRRRRRRRRRRRRRRRRCRRGMbFRRRRRRRRR>R=RbCGF
M,RRRRRRRRRRRRRRRRRRRRRRRRRo#HMRRRRRRRRRRR=#>RH,oM
RRRRRRRRRRRRRRRRRRRRRRRR0R#H$O	RRRRRRRRRR=>#O0H	
$,RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRRMRRoskN8RRRRRRRR>R=RkMoN2s8;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMMlFsNxDHC
;
R-R-Ro)CksDNRF"MsDlNH"xCRMVkOF0HMHRI0NERRH"#xsC_CR#"HkMb0R3
RMVkOF0HMFRMsDlNHRxC5R
RRsRVNRO0RRRRRRRRRRRRR:RRR)zh p1me_ 7zQh1t7h ;RRRRRRRRRRRR-RR-MRk#MHoCR8
RCRRGMbFRRRRRRRRRRRRRRRR:hRz)m 1p7e _t1Qh; 7R-R-RbCGFMMC0RR-4M,RFNslDCHx8R
RRHR#oRMRRRRRRRRRRRRRR:RRR71a_mzpt;QBR-R-Ro#HMHRL0R
RR0R#H$O	RRRRRRRRRRRRR:RRR71a_mzptRQB:'=RjR';RR--1O0H	L$RH50RsMFk8oHM2R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRR--k8#CRsVFRx#HHRMoF$MD
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0MM0RoskN8RRRR:RRRahqzp)qRRRR:V=RD0FN_NoksL8_H20#R-RR-kRoNRs8L#H0
RRRR0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sMMRFNslDCHxRs5VNRO0RRRRRRRRRR=>VOsN0R,
RRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=C>RGMbF,R
RRRRRRRRRRRRRRRRRRRRR#MHoRRRRRRRRR=RR>HR#o
M,RRRRRRRRRRRRRRRRRRRRR0R#H$O	RRRRRRRRRR=>#O0H	
$,RRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>-x#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=#>RH_xCs'C#EEHo,R
RRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRoRMk8NsRRRRRRRRRR=>MNoks;82
CRRMV8Rk0MOHRFMMlFsNxDHC
;
R-R-R0)Ck#sMRC0ERNOD#I#REEHORVXRN#DDR0HMFR
RVOkM0MHFRNBD#b#VRR5
RGRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RR-RR-DRVFHN0MboRF0HMRbHMkR0
RORRE	CO_sCsF:sRRmAmph qRR:=VNDF0E_OC_O	CFsssR2RRR--OOEC	FRVssRCs#Fs
RRRR0sCkRsMPHND8b_V#00NCR
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRaQh )t RR:=-MlHC'5GD,FIRDG'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERR:Q hatR ):G=R'oEHER;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRPHNsNCLDRoNsRRRRRRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RCRLoRHMRR--O#DN#
VbRRRRH5VRN'soDoCM0<ERRF4RssRVNHO0FIM_HE80Rd<RRRFsCFGbM0CM_8IH0<ERRRd
RRRRRFRRs'RGD0CVRG<R'osHER020MEC
RRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRRRRR&"qBp1u1w:RR"&R
RRRRRRwR"D0FNHRMobMFH0kRMlsLCR08CCCO08HRI0NERR8LNRMsNo
C"RRRRRRRR#CCPs$H0RsCsF
s;RRRRRCRs0MksRGH#;R
RRMRC8VRH;R
RR-R-RCBEOV	RF"sRX
"3RRRRNRso:0=RF4_jR,5GR''X2R;
RHRRVNR5sjo52RR='2X'RC0EMR
RRRRRskC0sHMR#RG;RRRRRRRRRRRRRRRRRRRRR-R-RRQV0sECC#RHRRNMXMRHRC0ERlMkL
CsRRRRR-R-RC1bODHNR#ONCR#,OOEC	FRVsDRHDNCoDkRMlsLC
RRRR#CDHOVRE	CO_sCsFNsRMR8
RRRRRM5N81R5az7_pQmtB _eB)amRs5NoCR5GMbFC_M0I0H8ER-48MFI0jFR2
22RRRRR=RRR''42ER0CRMRRRRRRRRRRRRRRRRRRRRR- -RGMbFCRM0HN#RD"DR4
"3RRRRRVRHRRFs5_0F#RDP5oNsR45-RI8FMR0F-NVsOF0HMH_I820E2R2
RRRRR/RR=jR''ER0CRMR-w-Rs0NOHRFMl0k#RRLCNRDD"Rj"F0sRERH#HM#RFN0RRlMkL3Cs
RRRRRRRRRHV5oNs52-4R'=R4R'20MECRRRRRRRRRR--wlsFR3"WRNiEMRR-Q   RN#0Ms8N8R
RRRRRRRRRskC0sMMRNRM;RRRRRRRRR-RR-6R(cHRLM$NsRRwu1MHoNMDHoNRMMhR5FN0RRlMkL2Cs
RRRRRRRR#CDCR
RRRRRRRRRskC0sJMRk0HC_MMN;R
RRRRRRMRC8VRH;R
RRRRRR-R-RCBEOV	RFHsRMMVHH
0$RRRRRDRC#RHVN5soCFGbM0CM_8IH0RE2=jR''ER0CRM
RRRRRsRRCs0kMFRb#M_HVR;RRRRRRRRRRRRRR-RR-FRu#HH0PHCRMMVHH
0$RRRRRDRC#RC
RRRRRsRRCs0kMCRMoM_HVR;RRRRRRRRRRRRRR-RR-CRhoHN0PHCRMMVHH
0$RRRRRMRC8VRH;R
RRRRR-O-RE	CORsVFR""j
RRRR#CDHFVRs1R5ap7_mBtQ_Be aRm)5oNsRG5CbCFMMI0_HE80-84RF0IMF2Rj2R2
RRRRR'=Rj0'RERCMRRRRRRRRRRRRRRRRRRRRR-RR-GR bCFMMH0R#DRNDjR""R
RRRRRHFVRs0R5FD_#PNR5s5oR-84RF0IMFVR-s0NOH_FMI0H8E222
RRRRRRRR'=Rj0'RERCMRRRRRRRRRRRRRRRRRRRRRR--wOsN0MHFRRH#NRDD"
j"RRRRRRRRHNVRsCo5GMbFC_M0I0H8E=2RR''jRC0EMR
RRRRRRRRRskC0sbMRFx#_C;sFRRRRRRRRRRRRR-R-RsZCFR
RRRRRRDRC#RC
RRRRRRRRR0sCkRsMM_CoxFCs;R
RRRRRRMRC8VRH;R
RRRRRCCD#
RRRRRRRRRHVN5soCFGbM0CM_8IH0RE2=jR''ER0CRM
RRRRRRRRR0sCkRsMb_F#8FCMsDlN;RRRRRRRR-RR-CR7MlFsNMDRkClLsHR5CRCCCCG0M88CR2Vb
RRRRRRRR#CDCR
RRRRRRRRRskC0sMMRC8o_CsMFl;ND
RRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RCRRD
#CRRRRRVRHRoNs5bCGFMMC0H_I820ER'=Rj0'RE
CMRRRRRRRRskC0sbMRFM#_FNslDR;RRRRRRRRRRRRR-h-RFNslDuRwRlMkL
CsRRRRRDRC#RC
RRRRRsRRCs0kMCRMoF_MsDlN;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8kRVMHO0FBMRD#N#V
b;
bRRsCFO8CksRCLsNM	_kClLs
R5RRRRNRsoRRRRRRRR:MRHRhRz)m 1p7e _FVDN
0;RRRR8FCMsDlNHRxC:MRHRmRAmqp h=R:RFVDN80_CsMFlHNDx
C;RRRROOEC	s_CsRFs:MRHRmRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRVOsN0RRRRRRR:kRF0hRz)m 1p7e _1zhQ th7R;
RCRRGMbFRRRRR:RRR0FkR)zh p1me_ 71hQt 
7;RRRR#MHoRRRRRRRR:kRF0aR17p_zmBtQ2#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=lR-H5MCN'soD,FIRoNs'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRPHNsNCLDR0Vb$RbRRRRRRRRR:NRPD_H8V0b#N;0C
LRRCMoH
RRRR0Vb$:bR=DRBNV##bNR5sRo,OOEC	s_Cs2Fs;R
RRHR#oRMR:0=RFj_G4s5Nos5NoH'Eo2E2;R
RRsRLC_N	MLklC5sR
RRRRNRRsRoRRRRRR=RR>sRNoR,
RRRRR0Vb$RbRRRRRRR=>V$b0bR,
RRRRRM8CFNslDCHxRR=>8FCMsDlNH,xC
RRRRVRRs0NORRRRR=RR>sRVN,O0
RRRRCRRGMbFRRRRR=RR>GRCb2FM;R
RCRM8bOsFCs8kCsRLC_N	MLklC
s;RRR
RFbsOkC8sLCRs	CN_lMkLRCs5R
RRsRNoRRRRRRRRRR:HRMRz h)1emp V7_D0FN;R
RRCR8MlFsNxDHCRR:HRMRApmm Rqh:V=RD0FN_M8CFNslDCHx;R
RREROC_O	CFsssRR:HRMRApmm Rqh:V=RD0FN_COEOC	_sssF;R
RRsRVNRO0RRRRRRR:FRk0z h)1emp k7_VCHG8R;R-4-RRI8FMR0F-NVsOF0HMH_I8
0ERRRRCFGbMRRRRRRR:kRF0hRz)m 1p7e _t1Qh; 7R-R-RbCGFMMC0H_I8-0E4FR8IFM0RRj
R#RRHRoMRRRRR:RRR0FkR71a_mzpt2QBR
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RH-lMNC5sDo'FRI,N'soD2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RPRRNNsHLRDCV$b0bRRRRRRRR:RRRDPNHV8_bN#00
C;RRRRPHNsNCLDRskVNRO0RRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH08ERF0IMF2Rj;-RR-MRk#MHoCV8Rs0NOH
FMRCRLo
HMRRRRV$b0b=R:RNBD#b#VRs5NoO,RE	CO_sCsF;s2
RRRRo#HM:RR=FR0_4Gj5oNs5oNs'oEHE;22
RRRRCLsNM	_kClLs
R5RRRRRsRNoRRRRRRRR>R=RoNs,R
RRRRRV$b0bRRRRRRR=V>Rbb0$,R
RRRRR8FCMsDlNHRxC=8>RCsMFlHNDx
C,RRRRRsRVNRO0RRRRR>R=RskVN,O0
RRRRCRRGMbFRRRRR=RR>GRCb2FM;R
RRsRVNRO058jRF0IMFVR-s0NOH_FMI0H8E:2R=VRkH8GCRV5ks0NO2R;
R8CMRFbsOkC8sLCRs	CN_lMkL;Cs
R
R-q-RsEH0lHC0OkRVMHO0F
M#RkRVMHO0F"MRN"L#RR5
RNRRs:oRR)zh p1me_ 7VNDF0R2RRRRRRRRRR-RR-DRVFHN0MboRF0HMRbHMkR0
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _FVDN50RN'sosoNMCR2;RR--skC#DR0
RoLCHRM
RHRRVNR5sDo'C0MoERR>j02RE
CMRRRRRCRs#0kDRRRRRRRRRRRR:0=RF4_jRs5No',RX;'2
RRRRsRRCD#k0NR5sEo'H2oERR:=';j'RRRRRRRRRR--#RC00REC#MHoR0LHRR0FbHF#0CHPRRRRRR
RRRRRskC0ssMRCD#k0R;
RCRRD
#CRRRRRCRs0MksRwhquR;
RCRRMH8RVR;
R8CMRMVkOF0HMNR"L;#"
R
R-Q-R R  (R6c"oMCNP0HCV"Rk0MOH
FMRkRVMHO0F"MR-5"R
RRRRoNsRz:Rh1) m pe7D_VF2N0RRRRRRRRRRRRRRRRRRRRRRRRR-R-RFVDNM0HoFRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0NR5sso'NCMo2R;R-s-RCD#k0R
RLHCoMR
RRVRHRs5NoC'DMEo0Rj>R2ER0CRM
RRRRR#sCkRD0RRRRRRRRR:RR=FR0_Rj45oNs,XR''
2;RRRRRCRs#0kDRs5NoH'EoRE2:M=RFs0RCD#k0NR5sEo'H2oE;RRRRR--HCMPs#0RHRoML
H0RRRRRCRs0MksR#sCk;D0
RRRR#CDCR
RRRRRskC0shMRq;wu
RRRR8CMR;HV
CRRMV8Rk0MOHRFM";-"
R
R-q-R808HH,FMR8N8#IR0FDRVFHN0MboRF0HMRlMkL#Cs
VRRk0MOHRFMNR885R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0RERRh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0ERRR:hzqa)Rqp:l=RNlGHkDl5'oEHEs,R'oEHER2;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRMOF#M0N08RN8NoksR8RRRRRR:RRRahqzp)qRR:=oskN8R;RRRRRR-RR-8RN8MRFCkRoNRs8L
H0RRRRPHNsNCLDRbDV0C$b,VRsbb0$CRR:PHND8b_V#00NCR;
RPRRNNsHLRDCVCbs#0kDRRRRRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLCsRVNDO0,sRVNsO0R:RRR1zhQ th7VR5s0NOH_FMI0H8E++4No88k8NsRI8FMR0FjR2;RR--VOsN0MHF#R
RRNRPsLHNDVCRs0NOOV,Rs0NO#RRR:hRz1hQt 57RVOsN0sD'NCMo2R;R-O-RF0M#NRM0NRM8#VEH0RC8PHNsNCLD#R
RRNRPsLHNDkCRsNVsOR0,ksDVNRO0:hRz1hQt 57RVOsN0MHF_8IH08ERF0IMF2Rj;R
RRNRPsLHNDkCRVOsN0RRRRRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH04E++8N8oskN8FR8IFM0R;j2
RRRRsPNHDNLCGRCbDFM,GRCbsFMR:RRRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2R-R-RbCGFMMC0R#
RPRRNNsHLRDCsbCGFRMRRRRRRRRRR1:RQ th7CR5GMbFC_M0I0H8EFR8IFM0R;j2R-R-R#sCkRD0CFGbM0CM
RRRRsPNHDNLCER#HGV0RRRRRRRRR:RRRt1QhR 75bCGFMMC0H_I8R0E8MFI0jFR2R;R-#-RE0HVRNVsOF0HMR#
RPRRNNsHLRDC#MHoRRRRRRRRRRRRR1:Raz7_pQmtBR;RRR--#MHoRRFV0RECFbk0kR0
RPRRNNsHLRDCD0CVsEHo0RRRRRRRRA:Rm mpqRh;RRRRRR--D0CVRRFssEHo0#RkCR8
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLC0R#H$O	RRRRRRRRR:RRR71a_mzpt;QBR-RR-FR]DR8#bOsCHF#HMFRVsFRskHM8MRo
RoLCHRMR-N-R808HH
FMRRRRH5VRVOsN0MHF_8IH0=ERRFjRs'RDDoCM0<ERRF(Rs'RsDoCM0<ERRR(20MEC
RRRRDRRV$b0b:CR=#RHGR;
RCRRD
#CRRRRRVRDbb0$C=R:RNOD#b#VR,5DRCOEOC	_sssF2R;
RRRRRbsV0C$bRR:=O#DN#RVb5Rs,OOEC	s_Cs2Fs;R
RRMRC8VRH;R
RRVRHRV5Dbb0$CRR=HR#GFssRV$b0b=CRRGH#2ER0CRM
RRRRRsVbCD#k0=R:R05FE#CsRR=>'2X';R
RRDRC#RHV5bDV0C$bRM=RNFMRsVRDbb0$CRR=JCkH0N_MMsRF
RRRRRRRRRRRs0Vb$RbC=NRMMsRFRbsV0C$bRJ=Rk0HC_MMN2R
RRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,4RRRRRsRFRV5Dbb0$CRR=b_F#HRMVNRM8s0Vb$RbC=CRMoM_HVR2
RRRRRRFs5bDV0C$bRM=RCHo_MNVRMs8RV$b0b=CRR#bF_VHM2ER0CRM
RRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-3.4,
RRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRDRC#RHV5bDV0C$bRb=RFH#_MFVRsVRsbb0$CRR=b_F#H2MVRC0EMRRR-G-RRH+RM=VRRVHM
RRRRVRRb#sCkRD0:b=RFH#_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRCHD#VDR5V$b0b=CRRoMC_VHMRRFss0Vb$RbC=CRMoM_HV02RERCMR-R-R-GRRVHMR-=RH
MVRRRRRbRVskC#D:0R=CRMoM_HVRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RCRRDV#HRV5Dbb0$CRR=M_CoxFCsR8NMRbsV0C$bRM=RCxo_C2sFRC0EMRRR---RjRR+-=jRR
-jRRRRRbRVskC#D:0R=CRMoC_xsbFVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRCCD#
RRRRDRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>0GF_jD452R,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRD0Vb$RbC:O=RD#N#V5bRD#sCH,xCRDVN#;C2RRRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRs#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4s
2,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRRbsV0C$bRR:=O#DN#RVb5Css#CHx,NRVD2#C;RRRRR--CFsssN#RDNsC8O$RE	COCR8
RRRRRCLsNM	_kClLs
R5RRRRRRRRNRsoRRRRRRRR=D>RsHC#x
C,RRRRRRRRV$b0bRRRRRRR=D>RV$b0b
C,RRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx
C,RRRRRRRRVOsN0RRRRRRR=k>RDNVsO
0,RRRRRRRRCFGbMRRRRRRR=C>RGMbFD
2;RRRRRsRVNDO0RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RR=FR50sEC#>R=R''j2R;
RRRRRNVsOR0D5NVsOF0HMH_I8+0ENo88k8NsRI8FMR0FNo88k8Ns2=R:RVkDs0NO;R
RRRRRLNsC	k_MlsLCRR5
RRRRRNRRsRoRRRRRR=RR>sRsCx#HCR,
RRRRRVRRbb0$RRRRR=RR>VRsbb0$CR,
RRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHCR,
RRRRRVRRs0NORRRRR=RR>sRkVOsN0R,
RRRRRCRRGMbFRRRRR=RR>GRCbsFM2R;
RRRRRNVsOR0sRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=R:R05FE#CsRR=>'2j';R
RRRRRVOsN05sRVOsN0MHF_8IH0NE+8k8oNRs88MFI0NFR8k8oN2s8RR:=kssVN;O0
RRRR#RRE0HVG=R:RG5CbDFM5bCGFMMC0H_I8-0E4&2RRbCGF2MDRC-RGMbFsR;
RRRRRRHV#VEH0<GRRs-VNDO0'oEHEER0CRM
RRRRRsRRCFGbMRRRRR:=CFGbMCs5GMbFC_M0I0H8E2-4RC&RGMbFsR;
RRRRRVRRs0NOORRRRR:=VOsN0
s;RRRRRRRRVOsN0R#RR=R:R05FE#CsRR=>'2j';RRR-N-R8x8RC
sFRRRRRRRRD0CVsEHo0=R:RDVN#
C;RRRRRRRR#O0H	R$RR=R:RRFs5NVsO20D;R
RRRRRCHD#VER#HGV0Rj<RRC0EMR
RRRRRRER#HGV0RRRR:-=RRH#EV;0G
RRRRRRRRNVsOR0#R:RR=ER#H_V0sEHo0VR5s0NOD0,RFM_H0CCosE5#HGV02
2;RRRRRRRRVOsN0RORR=R:RNVsO;0s
RRRRRRRRGsCbRFMR:RR=GRCbsFM5bCGFMMC0H_I8-0E4&2RRbCGF;Ms
RRRRRRRRVDC0osHE:0R=NRVD;#C
R--RRRRR#RR0	HO$RRRRR:=F5sRVOsN05DR0HF_Mo0CC#s5E0HVG82RF0IMF2Rj2R;
RRRRR#RR0	HO$RRRRR:=#DlNDNVsO50RVOsN0RD,0HF_Mo0CC#s5E0HVG;22
RRRRCRRDV#HRH#EVR0G=RRj0MEC
RRRRRRRRGsCbRFM:C=RGMbFDG5CbCFMMI0_HE80-R42&GRCbDFM;R
RRRRRR0R#H$O	RR:=';j'
RRRRRRRRRHVVOsN0>sRRNVsOR0D0MEC
RRRRRRRRVRRs0NOORRRRR:=VOsN0
s;RRRRRRRRRsRVN#O0RRRR:V=Rs0NODR;
RRRRRRRRRVDC0osHE:0R=NRVD;#C
RRRRRRRR#CDCR
RRRRRRRRRVOsN0RORR=R:RNVsO;0D
RRRRRRRRVRRs0NO#RRRRR:=VOsN0
s;RRRRRRRRRCRDVH0soRE0:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRCRRDV#HRH#EVR0G>sRVNsO0'oEHEER0CRM
RRRRRsRRCFGbMRRRRR:=CFGbMCD5GMbFC_M0I0H8E2-4RC&RGMbFDR;
RRRRRVRRs0NO#RRRRR:=5EF0CRs#='>Rj;'2R-RR-8RN8CRxsRF
RRRRRVRRs0NOORRRRR:=VOsN0
D;RRRRRRRRD0CVsEHo0=R:Rk0sCR;
RRRRR#RR0	HO$RRRRR:=F5sRVOsN0;s2
RRRRCRRDV#HRH#EVR0G>RRj0MEC
RRRRRRRRNVsOR0#R:RR=ER#H_V0sEHo0VR5s0NOs0,RFM_H0CCosE5#HGV02
2;RRRRRRRRVOsN0RORR=R:RNVsO;0D
RRRRRRRRGsCbRFMR:RR=GRCbDFM5bCGFMMC0H_I8-0E4&2RRbCGF;MD
RRRRRRRRVDC0osHE:0R=sR0k
C;-R-RRRRRR0R#H$O	RRRR:F=RsVR5s0NOs0R5FM_H0CCosE5#HGV02FR8IFM0R2j2;R
RRRRRR0R#H$O	RRRR:#=RlDNDVOsN0VR5s0NOs0,RFM_H0CCosE5#HGV02
2;RRRRRMRC8VRH;R
RRRRR-N-R8R8
RRRRRNVsOR0#5Rj2:V=Rs0NO#jR52sRFRH#0O;	$RRRRRR--m0sRE#CR0	HO$HRL0MRH00FREpCR1RA
RRRRRRHVD'5DEEHo2RR=s'5sEEHo2ER0CRM
RRRRRkRRVOsN0=R:RNVsOR0O+sRVN#O0;R
RRRRRRHR#oRMRRR:=D'5DEEHo2R;
RRRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-HR#oRM#NRsC8VHVCMsC0R
RRRRRRVRks0NORR:=VOsN0-ORRNVsO;0#RRRRR-R-RINDNR$#bHF#0CHPR#sCk
D0RRRRRRRRHDVRCsV0H0oERC0EMRRRRRRRRRRRRRRR-w-RHsokCkRF0ERIHROE#MHoRR0Fk
#CRRRRRRRRRHR#o:MR=5RDDH'Eo;E2
RRRRRRRR#CDCR
RRRRRRRRR#MHoRR:=s'5sEEHo2R;
RRRRRCRRMH8RVR;
RRRRR8CMR;HV
RRRRHRRVsRFRV5ks0NO2RR='Rj'0MEC
RRRRRRRRo#HM=R:R''j;RRRRRRRRRRRRRRRRRRRRR--Q   RcU6,3Rndb,RNosNsENbR
.3RRRRRMRC8VRH;R
RRRRR-M-RFNslDCHx
RRRRVRRb#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>kNVsO
0,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=s>RCFGbMR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRR#MHoRRRRRRRRR=RR>HR#o
M,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRH#0OR	$RRRRRRRR=#>R0	HO$R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRoRMk8NsRRRRRRRRRR=>No88k8Ns2R;
RCRRMH8RVR;
RsRRCs0kMbRVskC#D
0;RMRC8kRVMHO0FNMR8
8;
-RR-kR1LN0sOF0HMB,RN#DDR8"N8
"3RkRVMHO0F#MRksL0NRO05R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RR-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0oskN8RRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H0;-RR-kRMlsLCRRFVoskN8HRL0R#
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDMCRCRos:hRz)m 1p7e _FVDN50RsN'sM2oC;-RR-CRMoHN0PPCRCHs#FFMRV
RsRCRLo
HMRRRRMsCoRR:=-Rs;RRRRRRRRRRRRRRRRRRRRRRRR-s-RRR:=-Rs
RsRRCs0kM8RN8DR5RRRRRRRRR=RR>,RD
RRRRRRRRRRRRRRRRRsRRRRRRRRRRR=>MsCo,R
RRRRRRRRRRRRRRFRsk_M8#D0$C>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRkRoNRs8RRRRR>R=RNoks
8,RRRRRRRRRRRRRRRROOEC	s_CsRFs=O>RE	CO_sCsF
s,RRRRRRRRRRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx;C2
CRRMV8Rk0MOHRFM#0kLs0NO;R

RR--wNDF0oHMRHbFMl0RkHD0b
D$RkRVMHO0FlMRkHD0bRD$5R
RR,RDRRsRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0RERRh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0ERRR:hzqa)Rqp:l=RNlGHkDl5'oEHEs,R'oEHER2;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRMOF#M0N0kRlDk0oNRs8RRRRR:RRRahqzp)qRR:=oskN8R;RRRRRRRRRRR--oskN8HRL0R#
RPRRNNsHLRDCD0Vb$,bCRbsV0C$bRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDVCRb#sCkRD0RRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RRRRPHNsNCLDRNVsO,0DRNVsOR0sRRR:zQh1t7h Rs5VNHO0FIM_HE80RI8FMR0FjR2;RR--VOsN0MHF#R
RRNRPsLHNDsCRVOsN0RRRRRRRRRRR:hRz1hQt 57R55.*VOsN0MHF_8IH02E2+84RF0IMF2Rj;-RR-CRs#0kDRNVsOF0HMR
RRNRPsLHND#CRVOsN0RRRRRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH04E++Dlk0Noks88RF0IMF2Rj;-RR-CRs#0kDRNVsOF0HMR
RRNRPsLHND#CRE0HV$RRRRRRRRRRR:hRQa  t)R;RRRRR-8-RCsMFlRND#VEH0R
RRNRPsLHNDCCRGMbFDC,RGMbFsRRR:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2Rj;-RR-GRCbCFMM
0#RRRRPHNsNCLDRGsCbRFMRRRRRRRRRRR:1hQt 57RCFGbM0CM_8IH04E+RI8FMR0FjR2;RR--skC#DC0RGMbFC
M0RRRRPHNsNCLDR_Vb#MHoRRRRRRRRRRR:1_a7ztpmQRB;R-R-Ro#HMVRFR#sCk
D0RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RRNRPsLHND#CR0	HO$RRRRRRRRRRR:aR17p_zmBtQ;RRR-]-RF#D8RCbsOHH#FVMRFssRF8kMH
MoRCRLoRHMRR--l0kDH$bD
RRRRRHV5NVsOF0HMH_I8R0E=RRjFDsR'MDCoR0E<RR(FssR'MDCoR0E<2R(RC0EMR
RRRRRD0Vb$RbC:H=R#
G;RRRRCCD#
RRRRDRRV$b0b:CR=DRONV##bDR5,EROC_O	CFsss
2;RRRRRVRsbb0$C=R:RNOD#b#VR,5sRCOEOC	_sssF2R;
RCRRMH8RVR;
RHRRVDR5V$b0b=CRRGH#RRFss0Vb$RbC=#RHG02RE
CMRRRRRbRVskC#D:0R=FR50sEC#>R=R''X2R;
RCRRDV#HRD55V$b0b=CRRMMNRRFsD0Vb$RbC=kRJH_C0MRNMFRs
RRRRRRRRRsRRV$b0b=CRRMMNRRFss0Vb$RbC=kRJH_C0M2NM2ER0CRM
RRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-344,
RRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRDRC#RHV5D55V$b0b=CRR#bF_VHMRRFsD0Vb$RbC=CRMoM_HVN2RMR8
RRRRRRRRR5RRs0Vb$RbC=FRb#C_xsFFRsVRsbb0$CRR=M_CoxFCs2F2RsR
RRRRRRRRRRs55V$b0b=CRR#bF_VHMRRFss0Vb$RbC=CRMoM_HVN2RMR8
RRRRRRRRR5RRD0Vb$RbC=FRb#C_xsFFRsVRDbb0$CRR=M_CoxFCs2R220MECRRRR-j-RRH*RMRV
RRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-3d4,
RRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRDRC#RHV5bDV0C$bRb=RFH#_MFVRsVRsbb0$CRR=b_F#H
MVRRRRRRRRRFRRsVRDbb0$CRR=M_CoHRMVFssRV$b0b=CRRoMC_VHM2ER0CRMR-G-RRH*RM=VRRVHM
RRRRVRRb#sCkRD0:b=RFH#_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRR-R-RoVHkRsCFRk00REC#MHo
RRRRVRRbH_#o:MR=5RDDH'EoRE2GRFss'5sEEHo2R;RR-RR-HRVoCksR0FkRC0ERo#HMR
RRRRRVCbs#0kDRG5CbCFMMI0_HE802=R:R_Vb#MHo;R
RRDRC#RC
RRRRR_Vb#MHoRR:=D'5DEEHo2FRGs5RssH'Eo;E2RRRRRR--VkHosFCRk00RE#CRH
oMRRRRRsRDCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425D,R
RRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRDRRV$b0b:CR=DRONV##bDR5sHC#xRC,V#NDCR2;R-RR-sRCs#FsRsNDC$N8RCOEO8	C
RRRRsRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>0GF_js452R,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRs0Vb$RbC:O=RD#N#V5bRs#sCH,xCRDVN#;C2RRRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRLNsC	k_MlsLCRR5
RRRRRNRRsRoRRRRRR=RR>sRDCx#HCR,
RRRRRVRRbb0$RRRRR=RR>VRDbb0$CR,
RRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHCR,
RRRRRVRRs0NORRRRR=RR>sRVNDO0,R
RRRRRRGRCbRFMRRRRR>R=RbCGF2MD;R
RRRRRLNsC	k_MlsLCRR5
RRRRRNRRsRoRRRRRR=RR>sRsCx#HCR,
RRRRRVRRbb0$RRRRR=RR>VRsbb0$CR,
RRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHCR,
RRRRRVRRs0NORRRRR=RR>sRVNsO0,R
RRRRRRGRCbRFMRRRRR>R=RbCGF2Ms;R
RRRRRH5VRs0Vb$RbC=FRb#C_8MlFsNFDRsVRsbb0$CRR=M_Co8FCMsDlN2ER0CRM
RRRRR#RRE0HV$=R:RNVsOF0HMH_I8R0E-HRVMD8_ClV0F5#0VOsN0Rs,'24';R
RRRRRRsRVNsO0RR:=#VEH0C_DV50RVOsN0Rs,#VEH0;$2
RRRRCRRDV#HRV5Dbb0$CRR=b_F#8FCMsDlNRRFsD0Vb$RbC=CRMoC_8MlFsNRD20MEC
RRRRRRRRH#EVR0$:V=Rs0NOH_FMI0H8ERR-V8HM_VDC0#lF0s5VNDO0,4R''
2;RRRRRRRRVOsN0:DR=ER#H_V0D0CVRs5VNDO0,ER#H$V02R;
RRRRR#CDCR
RRRRRRER#H$V0RR:=jR;
RRRRR-RR-FRh00CRERN0NCR8MlFsNMDRkClLsRR*NCR8MlFsNMDRkClLs#RHRINDNR$#xFCs3R
RRRRRCRM8H
V;RRRRR-R-RDlk0DHb$R
RRRRR-N-R808RECCRGMbFC#M0
RRRRsRRCFGbM=R:R#sCHRxC5bCGF,MDRGsCb'FMDoCM0RE2+GRCbsFMR#-RE0HV$RR+4R;
RRRRRssVNRO0:V=Rs0NODRR*VOsN0Rs;RRRRR-RR-kRvDb0HD0$REVCRs0NOH
FMRRRRRVR#s0NORR:=sNVsO50RsNVsOE0'HRoE8MFI0RF
RRRRRRRRRRRRRRRRRRRRRsRRVOsN0H'Eo-ERRs5VNHO0FIM_HE80+l4+koD0k8Ns2
2;RRRRR0R#H$O	RR:=F5sRsNVsO50RsNVsOE0'H-oE5NVsOF0HMH_I8+0E4k+lDk0oN2s8
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2
2;RRRRR-R-RsMFlHNDxRC
RRRRRsVbCD#k0=R:RsMFlHNDx5CRVOsN0RRRRRRRR=RR>VR#s0NO,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFRRRRRRRRR>R=RGsCb,FM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRHR#oRMRRRRRRRRRRR=>V#b_H,oM
RRRRRRRRRRRRRRRRRRRRRRRRRRRR0R#H$O	RRRRRRRRRR=>#O0H	
$,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRRRRRRMRRoskN8RRRRRRRR>R=RDlk0Noks;82
RRRR8CMR;HV
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFRDlk0DHb$
;
RkRVMHO0F#MRE0Fs_P8HHR8C5R
RRGRD,GRsRz:Rht1Qh2 7
RRRR0sCkRsMzQh1t7h 
HRR#R
RR-R-RHaE##RHR#NRbHCON8DRH8PHCVsRF0sREVCRD0FNHRMobMFH0FRskM0HC
#3RRRR-w-RFNsRRk0sCMRk#MHoC88RH8PHCRs,"N#0o"C#RCMC80#RFRR=DEG'H
oERRRRO#FM00NMRN#0oRC#RRRRRRR:Q hatR ):D=RGH'Eo-ERR'sGEEHo;-RR-kRMlsLCRRFV#o0NCR#
RPRRNNsHLRDCb0NsHRNDRRRRRz:Rht1QhR 75'DGsoNMC
2;RRRRPHNsNCLDRRJRRRRRRRRRRRR:zQh1t7h R05#N#oCRI8FMR0Fj
2;RRRRPHNsNCLDRsbN0DHN_oNsDRR:1hQt 57RsEG'HRoE+RR.8MFI0jFR2R;
RPRRNNsHLRDCb0NsH_NDNRsoR1:RQ th7sR5GH'Eo+ERR8.RF0IMF2Rj;R
RLHCoMR
RRNRbsN0HD=R:R;DG
RRRRsVFRHHRM0R#N#oCRI8FMR0FjFRDFRb
RRRRRsbN0DHN_oNsD=R:R#sCHRxC5""jR1&RQ th7bR5NHs0NDD5GH'Eo8ERF0IMF2RH2R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsbN0DHN_oNsDC'DMEo02R;
RRRRRsbN0DHN_oNsRR:=b0NsH_NDNDsoR1-RQ th7"R5j&"RR2sG;R
RRRRRH5VRb0NsH_NDNRso5sbN0DHN_oNs'oEHE=2RR''42ER0CRMRRRRRRR--MNCo0CHP
RRRRRRRRHJ52=R:R''j;R
RRRRRCCD#
RRRRRRRRHJ52=R:R''4;R
RRRRRRNRbsN0HDDR5GH'EoHE+-N#0oRC#8MFI0DFRGH'EoHE+-N#0o-C#sEG'H2oER
:=RRRRRRRRRhRz1hQt 57Rb0NsH_NDN5sossG'NCMo2
2;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRR-0-RFNRl	0CREFCRkk0b0FRDFD	RHR	C00ENRRFV0RECkHM#o8MCR Q  HR8PCH83R
RRCRs0MksR#sCHRxC5RJ,DDG'C0MoE
2;RMRC8kRVMHO0F#MRE0Fs_P8HH;8C
R
R-4-R/VXRk0MOH3FMRCRhC88CRsVFRoNDF0sHE8lRCDPCFCblM
03RkRVMHO0FsMRCbOHsNFOD
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0kRoNRs8RRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0R#;RR--MLklCFsRVkRoNRs8L#H0
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RH-lMNC5sDo'FRI,N'soD2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=N'soEEHo;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RORRF0M#NRM08oHPk8NsRRRRR:RRRahqzp)qRR:=oskN8R;RR-RR-kRoNRs8L#H0
RRRRMVkOF0HMMRFCP8H$
R5RRRRRsRNoRR:zQh1t7h 2R
RRRRRskC0szMRht1Qh
 7RRRRHR#
RRRRRsPNHDNLCRRJRRR:zQh1t7h 5*5.N'soEEHo2R+48MFI0jFR2R;
RRRRRsPNHDNLCMRFCRR:zQh1t7h R'5JsoNMC
2;RRRRLHCoMR
RRRRRFRMCRRRRRRRRR=R:R05FE#CsRR=>'2j';R
RRRRRF5MCF'MCEEHo2=R:R''4;R
RRRRRJ=R:RF#Es80_H8PHCFR5MRC,N2so;RRRR-R-R#zMHCoM8HR8PCH8
RRRRsRRCs0kMCRs#CHxR,5JRoNs'MDCo+0E4
2;RRRRCRM8VOkM0MHFRCFM8$HP;R
RRNRPsLHNDVCRbb0$CRRRRRRRRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDCCRGMbFRRRRRRRRR1:RQ th7CR5GMbFC_M0I0H8ER-48MFI0jFR2R;RRR--CFGbM0CM#R
RRNRPsLHND8CRCsMFlV_FV0#CRh:Rq)azqspRNCMoR0jRF;R.
RRRRsPNHDNLCsRVNRO0RRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH08ERF0IMF2Rj;R
RRNRPsLHNDVCRs0NOoRRRRRRRRz:Rht1QhR 75NVsOF0HMH_I8+0E8oHPk8NsRI8FMR0Fj
2;RRRRPHNsNCLDRs#VNRO0RRRRR:RRR1zhQ th7VR5s0NOH_FMI0H8E++48oHPk8NsRI8FMR0FjR2;RR--skC#DV0Rs0NOH
FMRRRRPHNsNCLDRsVbCD#k0RRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RoLCHRMR-s-RCbOHsNFODR
RRbRV0C$bRR:=O#DN#5VbN,soRCOEOC	_sssF2R;
RORRD#N#OCN#RO:RNR#CV$b0bHCR#R
RRRRRIMECRGH#R
=>RRRRRRRRVCbs#0kDRR:=5EF0CRs#='>RX;'2
RRRRIRRERCMMRNM|kRJH_C0MRNM=R>
RRRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,R4
RRRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRERICbMRFH#_M|VRRoMC_VHMRR=>RRRRRRRR-4-R/VHM,CRs0MksRRj
RRRRRVRRb#sCkRD0:x=RCVsFbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRERICMMRCxo_CRsF|FRb#C_xs=FR>RRRRRRR-4-R/Rj
RRRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRRRRRR&)R" uBQ)qmBpw:RD0FNHRMouMFH0HR8PCH8RRL$xFCs"R
RRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRVCbs#0kDRR:=b_F#HVMVbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRCIEM0RFE#CsR
=>RRRRRRRRH5VRV$b0b=CRR#bF_M8CFNslDsRFR0Vb$RbC=CRMoC_8MlFsN
D2RRRRRRRRRMRN85R5NRso52-4RRFsN5so-2.2RR/='24'RC0EMR
RRRRRRRRR-4-R/M8CFNslDRR=HHMVM$H0,HRI00ERECCRGbOC0MHFRRFV.-**CFGbMN_L#RC
RRRRRRRRRsVbCD#k0=R:R#bF_VHMV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRRRRVCbs#0kDRG5CbCFMMI0_HE802=R:R_0FGRj45oNsRG5CbCFMMI0_HE802
2;RRRRRRRRCCD#
RRRRRRRRLRRs	CN_lMkLRCs5R
RRRRRRRRRRsRNoRRRRRRRR>R=RoNs,R
RRRRRRRRRRbRV0R$bRRRRR>R=R0Vb$,bC
RRRRRRRRRRRRM8CFNslDCHxRR=>8FCMsDlNH,xC
RRRRRRRRRRRRNVsOR0RRRRRRR=>VOsN0R,
RRRRRRRRRCRRGMbFRRRRR=RR>GRCb2FM;R
RRRRRRRRRVOsN0:oR=FR50sEC#>R=R''j2R;
RRRRRRRRRRHV50Vb$RbC=FRb#C_8MlFsNFDRsbRV0C$bRM=RC8o_CsMFl2NDRC0EMR
RRRRRRRRRR-R-RCaEROsCHFbsORNDFNVRRM8CFNslDkRMlsLCRRH#0H$bODND$CRxs
F,RRRRRRRRRRRR-C-RGbOC0FRVsIR0FbR#CNOHDNRO#RC#IOEHEsRNCsR0NCbb8CREs
C3RRRRRRRRRRRRH5VR0GF_jN45s5oR-242R'=R4R'20MEC
RRRRRRRRRRRRVRRs0NOoVR5s0NOoH'Eo8ERF0IMFHR8PNoks48+2=R:
RRRRRRRRRRRRRRRRNVsO50RVOsN0H'Eo4E-RI8FMR0FjR2;RRRRRR--1VEH0FR0R0MFRM8CFNslDR
RRRRRRRRRRRRR8FCMsFl_VCV#0=R:RR4;RRRRR-R-R8N8R04RFGRCbCFMMO0RFClbM0#NCR
RRRRRRRRRRDRC#RCRRRRRRRRRRRRRRRRRRRRRR-R-RoNs52-.R'=R4R'
RRRRRRRRRRRRRNVsOR0o5NVsO'0oEEHoRI8FMR0F8oHPk8Ns+R.2:R=
RRRRRRRRRRRRRVRRs0NORs5VN'O0EEHo-8.RF0IMF2Rj;RRRR-RR-ER1HRV00MFRF80RCsMFl
NDRRRRRRRRRRRRRCR8MlFs_VFV#RC0:.=R;RRRRRRR-N-R8.8RRR0FCFGbM0CMRlOFb#CMN
0CRRRRRRRRRRRRCRM8H
V;RRRRRRRRRDRC#RC
RRRRRRRRRVRRs0NOoVR5s0NOoH'Eo8ERF0IMFHR8PNoksR82:V=Rs0NO;R
RRRRRRRRRRCR8MlFs_VFV#RC0RRRRRRRRRRRRRRRRRRRRR:RR=;Rj
RRRRRRRRCRRMH8RVR;
RRRRRRRRRbCGFRMR:-=RRbCGF-MRR+dRRM8CF_slF#VVC
0;RRRRRRRRRVR#s0NORR:=F8MCHRP$5NVsO20o;R
RRRRRRRRR-M-RFNslDCHx
RRRRRRRRVRRb#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>#NVsO
0,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=C>RGMbF,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#RRHRoMRRRRRRRRR>R=RoNs5bCGFMMC0H_I820E,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#RR0	HO$RRRRRRRR>R=R''4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRkMoNRs8RRRRRRRR=8>RHkPoN2s8;R
RRRRRRMRC8VRH;R
RRMRC8NRO#OCRD#N#OCN#;R
RRCRs0MksRsVbCD#k0R;
R8CMRMVkOF0HMCRsOsHbFDON;R

RR--VNDF0oHMRHbFM80RH#PHH
FMRkRVMHO0F8MRH8PHC
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0RRRRR-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0oskN8RRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H0;-RR-kRMlsLCRRFVoskN8HRL0R#
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRFROMN#0MV0Rs0NOH_FMI0H8ERRR:qRhaqz)p=R:RH-lMDC5'IDF,'RsD2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0RERRh:Rq)azq:pR=NRlGkHll'5DEEHo,'RsEEHo2R;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRO#FM00NMRP8HoskN8RRRRRRRRRR:hzqa)Rqp:o=Rk8Ns;-RR-HR8PHH#FoMRk8NsR0LH#R
RRNRPsLHNDDCRV$b0bRC,s0Vb$RbC:NRPD_H8V0b#N;0C
RRRRsPNHDNLCbRVskC#DR0RRRRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RPRRNNsHLRDCksDVN,O0RVkss0NORz:Rht1QhR 75NVsOF0HMH_I8R0E8MFI0jFR2R;
RPRRNNsHLRDCVOsN0RDRRRRRRRRRRz:Rht1QhR 75*5.5NVsOF0HMH_I8+0E8oHPk8Ns22+4RI8FMR0FjR2;RR--D0CV
RRRRsPNHDNLCsRVNsO0RRRRRRRRR:RRR1zhQ th7VR5s0NOH_FMI0H8EH+8PNoks88RF0IMF2Rj;-RR-HRso
E0RRRRPHNsNCLDRssVNRO0RRRRRRRRRRR:zQh1t7h Rs5VNDO0'MsNo;C2RRRR-s-RCD#k0sRVNHO0FRM
RPRRNNsHLRDC#NVsOR0RRRRRRRRRRz:Rht1QhR 75NVsOF0HMH_I8+0E4H+8PNoks88RF0IMF2Rj;-RR-CRs#0kDRNVsOF0HMR
RRNRPsLHNDCCRGMbFDC,RGMbFsRRR:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2Rj;-RR-GRCbCFMM
0#RRRRPHNsNCLDRGsCbRFMRRRRRRRRRRR:1hQt 57RCFGbM0CM_8IH04E+RI8FMR0FjR2;RR--skC#DC0RGMbFC
M0RRRRPHNsNCLDR_Vb#MHo,0R#H$O	RRR:1_a7ztpmQRB;RRRRR-RR-HR#oFMRVCRs#0kD
RRRRsPNHDNLCER#H$V0,ER#HGV0R:RRRaQh )t ;RRRRRRRRRRR-8-RCsMFlRNDMLklC#sRE0HV
RRRRsPNHDNLCsRDCx#HCs,RsHC#x:CRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RoLCHRMR-8-RH8PHCR
RRVRHRs5VNHO0FIM_HE80Rj=RRRFsDC'DMEo0R(<RRRFssC'DMEo0R(<R2ER0CRM
RRRRRbDV0C$bRR:=H;#G
RRRR#CDCR
RRRRRD0Vb$RbC:O=RD#N#V5bRDO,RE	CO_sCsF;s2
RRRRsRRV$b0b:CR=DRONV##bsR5,EROC_O	CFsss
2;RRRRCRM8H
V;RRRRO#DN##ONCRR:OCN#RbsV0C$bR
H#RRRRRERICHMR#=GR>R
RRRRRRbRVskC#D:0R=FR50sEC#>R=R''X2R;
RRRRRCIEMNRMMRR|JCkH0N_MM>R=
RRRRRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-344,
RRRRRRRRsVbCD#k0=R:RNJMMRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRIMECR#bF_VHMRM|RCHo_M=VR>R
RRRRRRVRHRbDV0C$bRb=RFH#_MFVRsVRDbb0$CRR=M_CoHRMVRR--HRMV/MRHVR
RRRRRRRRRFDsRV$b0b=CRRHJkCM0_NFMRsVRDbb0$CRR=MRNM0MEC
RRRRRRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,Rc
RRRRRRRRRsVbCD#k0=R:RNJMMRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRR-G-RRH/RM=VRRRj
RRRRRRRRRsVbCD#k0=R:RsxCFRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRRbRV_o#HM=R:RDD5'oEHEG2RFssR5Es'H2oE;RRRRRRRRR--#MHo
RRRRRRRRVRRb#sCkRD05sVbCD#k0H'EoRE2:V=RbH_#oRM;RR--#MHo
RRRRRRRR8CMR;HV
RRRRIRRERCMb_F#xFCsRM|RCxo_CRsF=R>
RRRRRHRRVVRDbb0$CRR=b_F#xFCsRRFsD0Vb$RbC=CRMoC_xsRFRRRRRR-RR-RRj/
RjRRRRRRRRRsRFRbDV0C$bRJ=Rk0HC_MMNRRFsD0Vb$RbC=NRMMER0CRM
RRRRRRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-3c4,
RRRRRRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRDRC#RC
RRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRRRRRR&7R"Q7eQ w:RD0FNHRMouMFH0HR8PCH8RRL$xFCs"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRR-Q-RMMVHH,0$RV8CHRMCH(MR64c-g-U6(
3.RRRRRRRRRbRVskC#D:0R=FRb#M_HVRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRRRRR_Vb#MHoRR:=D'5DEEHo2FRGs5RssH'Eo;E2RRRRRRRR-#-RH
oMRRRRRRRRRbRVskC#D50RVCbs#0kD'oEHE:2R=bRV_o#HMR;R-#-RH
oMRRRRRRRRCRM8H
V;RRRRRERICFMR0sEC#>R=
RRRRRRRRNOD#N#O#RC.:NRO#DCRV$b0bHCR#R
RRRRRRRRRIMECRGH#R
=>RRRRRRRRRRRRVCbs#0kDRR:=5EF0CRs#='>RX;'2
RRRRRRRRIRRERCMMRNM|kRJH_C0MRNM=R>
RRRRRRRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,R4
RRRRRRRRRVRRb#sCkRD0:J=RMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRRERICbMRFH#_M|VRRoMC_VHMRR=>RRRR-H-RM/VRR=GRRVHM
RRRRRRRRRRRRsVbCD#k0=R:R#bF_VHMV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRRRRRV#b_HRoM:D=R5ED'H2oERsGFRss5'oEHER2;RRRRR-RR-HR#oRM
RRRRRRRRRVRRb#sCk5D0CFGbM0CM_8IH0RE2:V=RbH_#o
M;RRRRRRRRRERICbMRFx#_CRsF|CRMoC_xs=FR>RRR-j-RRX/RRj=R
RRRRRRRRRRRRsVbCD#k0=R:RsxCFRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRRRRRbRV_o#HM=R:RDD5'oEHEG2RFssR5Es'H2oE;RRRRRRRRR--#MHo
RRRRRRRRRRRRsVbCD#k0G5CbCFMMI0_HE802=R:R_Vb#MHo;R
RRRRRRRRRIMECREF0CRs#=R>
RRRRRRRRRVRRbH_#o:MR=5RDDH'EoRE2GRFss'5sEEHo2R;RRRRRR-R-Ro#HMR
RRRRRRRRRRsRDCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRRRRRRRRRbDV0C$bRR:=O#DN#RVb5CDs#CHx,NRVD2#C;RRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRRRRRRsRsCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425s,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRRRRRRRRRbsV0C$bRR:=O#DN#RVb5Css#CHx,NRVD2#C;RRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRRRRRRsRLC_N	MLklC5sR
RRRRRRRRRRRRNRRsRoRRRRRR=RR>sRDCx#HCR,
RRRRRRRRRRRRR0Vb$RbRRRRRRR=>D0Vb$,bC
RRRRRRRRRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRNVsOR0RRRRRRR=>ksDVN,O0
RRRRRRRRRRRRCRRGMbFRRRRR=RR>GRCbDFM2R;
RRRRRRRRR-RR-HRsoRE0#CH8
RRRRRRRRRRRRCLsNM	_kClLs
R5RRRRRRRRRRRRRsRNoRRRRRRRR>R=RCss#CHx,R
RRRRRRRRRRRRRV$b0bRRRRRRR=s>RV$b0b
C,RRRRRRRRRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRVOsN0RRRRRRR=k>RsNVsO
0,RRRRRRRRRRRRRGRCbRFMRRRRR>R=RbCGF2Ms;R
RRRRRRRRRR-R-RlBFbCk0RC0ERbCGFMMC0R
RRRRRRRRRRCRsGMbFRR:=sHC#x5CRCFGbMRD,sbCGFDM'C0MoE-2RRbCGFRMs-;R.
RRRRRRRRRRRRRHV5bsV0C$bRb=RF8#_CsMFlRNDFssRV$b0b=CRRoMC_M8CFNslD02RE
CMRRRRRRRRRRRRR-R-RR7F0REC#VEH0oHMRsECCFRM0VRN03CsRERaNI0RNI$RCNREPNCRRN#lDsDC
RRRRRRRRRRRR-RR-ER#HCV0sN,RMM8RCRC8NlR#NCDDsHR8PCH8sL,RCkON#0CRE0CRFRb
RRRRRRRRRRRRRR--LRH0H0MRE8CRH#PHFIsRHRDDNNDI$L#RCRRN"34"
RRRRRRRRRRRR#RRE0HV$=R:RNVsOF0HMH_I8R0E-HRVMD8_ClV0F5#0kssVN,O0R''42R;
RRRRRRRRRRRRRVkss0NORR:=#VEH0C_DV50RkssVN,O0RH#EV20$;R
RRRRRRRRRRRRRsbCGF:MR=CRsGMbFR#+RE0HV$R;
RRRRRRRRRCRRMH8RVR;
RRRRRRRRRVRRs0NOs=R:R05FE#CsRR=>'2j';R
RRRRRRRRRRsRVNsO0Rs5VNHO0FIM_HE80+P8HoskN8FR8IFM0RP8HoskN8:2R=sRkVOsN0R;
RRRRRRRRRHRRVDR5V$b0b=CRR#bF_M8CFNslDsRFRbDV0C$bRM=RC8o_CsMFl2NDRC0EMR
RRRRRRRRRRRRR#VEH0:GR=sRVNHO0FIM_HE80RV-RH_M8D0CVl0F#5VkDs0NO,4R''
2;RRRRRRRRRRRRRDRkVOsN0=R:RH#EVD0_CRV05VkDs0NO,ER#HGV02R;
RRRRRRRRRRRRRGsCbRFM:s=RCFGbMRR-#VEH0
G;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRVOsN0RDR:5=RFC0Es=#R>jR''
2;RRRRRRRRRRRRVOsN05DRVOsN0ED'HRoE8MFI0VFRs0NODH'EoVE-s0NOH_FMI0H8E:2R=DRkVOsN0R;
RRRRRRRRR-RR-HR8PCH8
RRRRRRRRRRRRssVNRO0:#=RE0Fs_P8HHR8C5NVsO,0DRNVsO20s;RRRRRRRRR--kHM#o8MCRP8HH
8CRRRRRRRRRRRR#NVsO:0R=VRss0NORV5#s0NO'MsNo;C2RRRRR-RR-FRDIRCsL#H0
RRRRRRRRRRRRH#0OR	$:'=R4
';RRRRRRRRRRRR-M-RFNslDCHx
RRRRRRRRRRRRsVbCD#k0=R:RsMFlHNDx5CRVOsN0RRRRRRRR=RR>VR#s0NO,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=s>RCFGbMR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRHR#oRMRRRRRRRRRRR=>V#b_H,oM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#O0H	R$RRRRRR=RR>0R#H$O	,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRRoskN8RRRRRRRR>R=RP8HoskN8
2;RRRRRRRRCRM8OCN#RNOD#N#O#;C.
RRRR8CMR#ONCDRONO##N;#C
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFRP8HH;8C
R
R-8-RH#PHHRFMLN$RRIbFCFsRV
R.RkRVMHO0F8MRH8PHCbL$.
R5RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0RRRRR-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0Mo0Rk8NsRRRRR:RRRahqzp)qRRRR:V=RD0FN_NoksL8_H;0#R-R-RlMkLRCsFoVRk8NsR0LH#R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80R:RRRahqzp)qRR:=-MlHC'5DD,FIRDs'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERRR:qRhaqz)p=R:RGlNHllk5ED'H,oEREs'H2oE;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RPRRNNsHLRDCD0Vb$,bCRbsV0C$bRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDVCRb#sCkRD0RRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RRRRPHNsNCLDRVkDs0NO,sRkVOsN0RR:zQh1t7h Rs5VNHO0FIM_HE80RI8FMR0Fj
2;RRRRPHNsNCLDRbCGF,MDRbCGFRMsRRR:1hQt C75GMbFC_M0I0H8ER-48MFI0jFR2R;R-C-RGMbFC#M0
RRRRsPNHDNLCCRsGMbFRRRRRRRRR:RRRt1Qh5 7CFGbM0CM_8IH08ERF0IMF2Rj;-RR-CRs#0kDRbCGFMMC0R
RRNRPsLHNDVCRbH_#oRMRRRRRRRRR:aR17p_zmBtQ;RRRRRRR-#-RHRoMFsVRCD#k0R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RCRLoRHMRR--8HHP#MHFL.$b
RRRRRHV5NVsOF0HMH_I8R0E=RRjFDsR'MDCoR0E<RR(FssR'MDCoR0E<2R(RC0EMR
RRRRRD0Vb$RbC:H=R#
G;RRRRCCD#
RRRRDRRV$b0b:CR=DRONV##bDR5,EROC_O	CFsss
2;RRRRRVRsbb0$C=R:RNOD#b#VR,5sRCOEOC	_sssF2R;
RCRRMH8RVR;
RORRD#N#OCN#RO:RNR#Cs0Vb$RbCHR#
RRRRRCIEM#RHG>R=
RRRRRRRRsVbCD#k0=R:R05FE#CsRR=>'2X';R
RRRRRIMECRMMNRJ|Rk0HC_MMNR
=>RRRRRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,4RRRRRRRRVCbs#0kDRR:=JMMNV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRIRRERCMb_F#HRMV|CRMoM_HV>R=
RRRRRRRRRHVD0Vb$RbC=FRb#M_HVsRFRbDV0C$bRM=RCHo_M0VRERCMRRRRRR--HRMV/MRHVR
RRRRRRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,cRRRRRRRRRbRVskC#D:0R=MRJNbMVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--GRR/HRMV=
RjRRRRRRRRRbRVskC#D:0R=CRxsbFVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRVRRbH_#o:MR=5RDDH'EoRE2GRFss'5sEEHo2R;RRRRRR-R-Ro#HMR
RRRRRRRRRVCbs#0kDRb5VskC#DE0'H2oERR:=V#b_H;oMR-R-Ro#HMR
RRRRRRMRC8VRH;R
RRRRRIMECR#bF_sxCFRR|M_CoxFCsR
=>RRRRRRRRHDVRV$b0b=CRR#bF_sxCFsRFRbDV0C$bRM=RCxo_CRsF0MECRRRR-j-RRj/R
RRRRRRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,Rc
RRRRRRRRRsVbCD#k0=R:RNJMMRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRCCD#
RRRRRRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRRRRRRRRR&"e7QQA7 Y:u.RFwDNM0HoFRuHRM08HHP8LCR$CRxs
F"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRR-R-RVQMH0MH$8,RCMVHCMRHRc(6-U4g63-(.R
RRRRRRRRRVCbs#0kDRR:=b_F#HVMVbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRVRRbH_#o:MR=5RDDH'EoRE2GRFss'5sEEHo2R;RRRRRR-R-Ro#HMR
RRRRRRRRRVCbs#0kDRb5VskC#DE0'H2oERR:=V#b_H;oMR-R-Ro#HMR
RRRRRRMRC8VRH;R
RRRRRIMECREF0CRs#=R>
RRRRRORRD#N#OCN#.RR:OCN#RbDV0C$bR
H#RRRRRRRRRERICHMR#=GR>R
RRRRRRRRRRbRVskC#D:0R=FR50sEC#>R=R''X2R;
RRRRRRRRRCIEMNRMMRR|JCkH0N_MM>R=
RRRRRRRRRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-344,
RRRRRRRRRRRRsVbCD#k0=R:RNJMMRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRRRRIMECR#bF_VHMRM|RCHo_M=VR>RRRR-R-RVHMRG/RRH=RMRV
RRRRRRRRRVRRb#sCkRD0:b=RFH#_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRRRRRbRV_o#HM=R:RDD5'oEHEG2RFssR5Es'H2oE;RRRRRRRRR--#MHo
RRRRRRRRRRRRsVbCD#k0CR5GMbFC_M0I0H8E:2R=bRV_o#HMR;R-#-RH
oMRRRRRRRRRERICbMRFx#_CRsF|CRMoC_xs=FR>RRR-j-RRX/RRj=R
RRRRRRRRRRRRsVbCD#k0=R:RsxCFRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRRRRRRRRRbRV_o#HM=R:RDD5'oEHEG2RFssR5Es'H2oE;RRRRRRRRR--#MHo
RRRRRRRRRRRRsVbCD#k0CR5GMbFC_M0I0H8E:2R=bRV_o#HMR;R-#-RH
oMRRRRRRRRRERICFMR0sEC#>R=
RRRRRRRRRRRR_Vb#MHoRR:=D'5DEEHo2FRGs5RssH'Eo;E2RRRRRRRR-#-RH
oMRRRRRRRRRRRRD#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4D
2,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRRRRRRDRRV$b0b:CR=DRONV##bDR5sHC#xRC,V#NDCR2;RR--CFsssN#RDNsC8O$RE	COCR8
RRRRRRRRRsRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>0GF_js452R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNH_xCH=MR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRRRRRRVRsbb0$C=R:RNOD#b#VRs5sCx#HCV,RNCD#2R;R-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRRRRRRsRLC_N	MLklC5sR
RRRRRRRRRRRRNRRsRoRRRRRR=RR>sRDCx#HCR,
RRRRRRRRRRRRR0Vb$RbRRRRRRR=>D0Vb$,bC
RRRRRRRRRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRNVsOR0RRRRRRR=>ksDVN,O0
RRRRRRRRRRRRCRRGMbFRRRRR=RR>GRCbDFM2R;
RRRRRRRRR-RR-HRsoRE0#CH8
RRRRRRRRRRRRCLsNM	_kClLs
R5RRRRRRRRRRRRRsRNoRRRRRRRR>R=RCss#CHx,R
RRRRRRRRRRRRRV$b0bRRRRRRR=s>RV$b0b
C,RRRRRRRRRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRVOsN0RRRRRRR=k>RsNVsO
0,RRRRRRRRRRRRRGRCbRFMRRRRR>R=RbCGF2Ms;R
RRRRRRRRRR#RN#0CsRs5FRs5kVOsN0VR5s0NOH_FMI0H8ER-48MFI0jFR2=2RR''j2R
RRRRRRRRRRRRRsFCbsw0Rpamq_ht  B)Q_tui'#HM0ONMCN_MlRC
RRRRRRRRRRRRR"&R7QQe7Y AuR.:"R
RRRRRRRRRRRRR&7R"H8PHCbL$.NROD8DCR0IHERRNMRFMbCFIsVRFRF0IRP8HHs#F"R
RRRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRRRRsbCGF:MR=CR5GMbFDG5CbDFM'oEHEC2&GMbFDR2
RRRRRRRRRRRRRRRRRRRRR5-RCFGbMCs5GMbFsH'Eo&E2CFGbMRs2-;R4
RRRRRRRRRRRRR--MlFsNxDHCR
RRRRRRRRRRbRVskC#D:0R=FRMsDlNHRxC5NVsOR0RRRRRRRRR=k>RDNVsO
0,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFRRRRRRRRR>R=RGsCb,FM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#MHoRRRRRRRRR=RR>bRV_o#HMR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR0R#H$O	RRRRRRRRRR=>',4'
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRoRMk8NsRRRRRRRRRR=>j
2;RRRRRRRRCRM8OCN#RNOD#N#O#;C.
RRRR8CMR#ONCDRONO##N;#C
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFRP8HHL8C$;b.
R
R-v-RkHD0bRD$NkOOlNkD0RCRskC#D=0RRsD*RO+R
VRRk0MOHRFMlRNO5R
RR,RDRRs,ORRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qR
:=RRRRRlR-HRMC5MlHC'5DD,FIRDs'F,I2RDO'F;I2R-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qR
:=RRRRRNRlGkHlllR5NlGHkDl5'oEHEs,R'oEHER2,OH'Eo;E2R-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHNDDCRV$b0bRC,s0Vb$,bCRbOV0C$bRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDVCRb#sCkRD0RRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLCsRVNDO0,sRVNsO0RRRRRRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH08ERF0IMF2Rj;-RR-sRVNHO0F
M#RRRRPHNsNCLDRNVsOR0GRRRRRRRRRRRRRRRRR:RRR1zhQ th7VR5s0NOH_FMI0H8Ek+oNRs88MFI0jFR2R;
RPRRNNsHLRDCVOsN0RO,VOsN0R#RRRRRRRRRRRR:zQh1t7h Rs5VNHO0FIM_HE80+o4+k8NsRI8FMR0Fj
2;RRRRPHNsNCLDRssVNRO0RRRRRRRRRRRRRRRRR:RRR1zhQ th75R5.V*5s0NOH_FMI0H8E+224FR8IFM0R;j2R-R-R#sCkRD0VOsN0MHF
RRRRsPNHDNLCVR#s0NO,VRks0NORRRRRRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH04E++Noks88RF0IMF2Rj;-RR-CRs#0kDRNVsOF0HMR
RRNRPsLHNDCCRGMbFDC,RGMbFsC,RGMbFORRRR1:RQ th7CR5GMbFC_M0I0H8ER-48MFI0jFR2R;R-C-RGMbFC#M0
RRRRsPNHDNLCCRsGMbF,CRsGMbF.RRRRRRRRRRR:QR1t7h RG5CbCFMMI0_HE80+84RF0IMF2Rj;-RR-CRs#0kDRbCGFMMC0R
RRNRPsLHND#CRE0HV$RRRRRRRRRRRRRRRRRRRRQ:Rhta  R);RRRRRR--8FCMsDlNRH#EVR0
RPRRNNsHLRDC#VEH0RGRRRRRRRRRRRRRRRRRRRR:1hQt 57RsbCGFsM'NCMo2R;R-#-RE0HVRNVsOF0HMR#
RPRRNNsHLRDCV#b_HRoMRRRRRRRRRRRRRRRRRRR:1_a7ztpmQRB;RR--#MHoRRFVskC#DR0
RPRRNNsHLRDCD#sCH,xCRCss#CHxRRRRRRRRRRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RRNRPsLHNDOCRsHC#xRCRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0-ERRNoks;82
RRRRsPNHDNLCCRDVH0soRE0RRRRRRRRRRRRRRRR:mRAmqp hR;RR-RR-CRDVF0RsHRsoRE0k8#C
RRRRsPNHDNLC0R#H$O	RRRRRRRRRRRRRRRRRRRR:aR17p_zmBtQ;-RR-FR]DR8#bOsCHF#HMFRVsFRskHM8MRo
RPRRNNsHLRDC#s0N0GH8:MRH0CCosR;
RoLCHRMR-l-RkHD0b
D$RRRRH5VRVOsN0MHF_8IH0=ERRFjRs'RDDoCM0<ERRF(Rs'RsDoCM0<ERRF(Rs'RODoCM0<ERRR(20MEC
RRRRDRRV$b0b:CR=#RHGR;
RCRRD
#CRRRRRVRDbb0$C=R:RNOD#b#VR,5DRCOEOC	_sssF2R;
RRRRRbsV0C$bRR:=O#DN#RVb5Rs,OOEC	s_Cs2Fs;R
RRRRRO0Vb$RbC:O=RD#N#V5bROO,RE	CO_sCsF;s2
RRRR8CMR;HV
RRRRRHV5bDV0C$bRH=R#FGRsVRsbb0$CRR=HR#GFOsRV$b0b=CRRGH#2ER0CRM
RRRRRsVbCD#k0=R:R05FE#CsRR=>'2X';R
RRDRC#RHV5bDV0C$bRM=RNFMRsVRDbb0$CRR=JCkH0N_MMsRF
RRRRRRRRRRRs0Vb$RbC=NRMMsRFRbsV0C$bRJ=Rk0HC_MMNR
FsRRRRRRRRRORRV$b0b=CRRMMNRRFsO0Vb$RbC=kRJH_C0M2NMRC0EMR
RRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,4RRRRRbRVskC#D:0R=MRJNbMVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRR#CDH5VR5V5Dbb0$CRR=b_F#HRMVFDsRV$b0b=CRRoMC_VHM2MRN8R
RRRRRRRRRRsR5V$b0b=CRR#bF_sxCFsRFRbsV0C$bRM=RCxo_C2sF2sRF
RRRRRRRRRRR5V5sbb0$CRR=b_F#HRMVFssRV$b0b=CRRoMC_VHM2MRN8R
RRRRRRRRRRDR5V$b0b=CRR#bF_sxCFsRFRbDV0C$bRM=RCxo_C2sF202RERCMRR--jRR*H
MVRRRRR-R-R0)CkRsMJCkH0qRhhQ,R (  64c-g-U6(,34dR
RRRRRVCbs#0kDRR:=JMMNV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RCRRDV#HRV5Dbb0$CRR=b_F#HRMVFssRV$b0b=CRR#bF_VHM
RRRRRRRRRRRFDsRV$b0b=CRRoMC_VHMRRFss0Vb$RbC=CRMoM_HV-RR-RRG*MRHVRR=H
MVRRRRRRRRRFRRsVRObb0$CRR=M_CoHRMVFOsRV$b0b=CRR#bF_VHM2ER0CRMR-G-RRH+RM=VRRVHM
RRRRVRRb#sCkRD0:b=RFH#_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRR-R-RoVHkRsCFRk00REC#MHo
RRRRVRRb#sCkRD05bCGFMMC0H_I820ERR:=D'5DEEHo2FRGs5RssH'Eo;E2
RRRR#CDCR
RRRRRV#b_HRoM:D=R5ED'H2oERsGFRss5'oEHER2;RR--VkHosFCRk00RE#CRH
oMRRRRRsRDCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425D,R
RRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRDRRV$b0b:CR=DRONV##bDR5sHC#xRC,V#NDCR2;RRRRR-RR-sRCs#FsRsNDC$N8RCOEO8	C
RRRRsRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>0GF_js452R,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRs0Vb$RbC:O=RD#N#V5bRs#sCH,xCRDVN#;C2RRRRRRRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRO#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4O
2,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>OR-sHC#xDC'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRORRV$b0b:CR=DRONV##bOR5sHC#xRC,V#NDCR2;RRRRR-RR-sRCs#FsRsNDC$N8RCOEO8	C
RRRRLRRs	CN_lMkLRCs5R
RRRRRRsRNoRRRRRRRR>R=RCDs#CHx,R
RRRRRRbRV0R$bRRRRR>R=RbDV0C$b,R
RRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRsRVNRO0RRRRR>R=RNVsO,0D
RRRRRRRRbCGFRMRRRRRRR=>CFGbM;D2
RRRRLRRs	CN_lMkLRCs5R
RRRRRRsRNoRRRRRRRR>R=RCss#CHx,R
RRRRRRbRV0R$bRRRRR>R=RbsV0C$b,R
RRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRsRVNRO0RRRRR>R=RNVsO,0s
RRRRRRRRbCGFRMRRRRRRR=>CFGbM;s2
RRRRLRRs	CN_lMkLRCs5R
RRRRRRsRNoRRRRRRRR>R=RCOs#CHx,R
RRRRRRbRV0R$bRRRRR>R=RbOV0C$b,R
RRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRsRVNRO0RRRRR>R=RNVsO,0G
RRRRRRRRbCGFRMRRRRRRR=>CFGbM;O2
RRRRHRRVsR5V$b0b=CRR#bF_M8CFNslDsRFRbsV0C$bRM=RC8o_CsMFl2NDRC0EMR
RRRRRRER#H$V0RR:=VOsN0MHF_8IH0-ERRMVH8C_DVF0l#V05s0NOs',R4;'2
RRRRRRRRNVsOR0s:#=RE0HV_VDC0VR5s0NOs#,RE0HV$
2;RRRRRDRC#RHV5bDV0C$bRb=RF8#_CsMFlRNDFDsRV$b0b=CRRoMC_M8CFNslD02RE
CMRRRRRRRR#VEH0:$R=sRVNHO0FIM_HE80RV-RH_M8D0CVl0F#5NVsO,0DR''42R;
RRRRRVRRs0NOD=R:RH#EVD0_CRV05NVsO,0DRH#EV20$;R
RRRRRCCD#
RRRRRRRRH#EVR0$:j=R;R
RRRRRR-R-R0hFCER0NN0RRM8CFNslDkRMlsLCRN*RRM8CFNslDkRMlsLCRRH#NNDI$x#RC3sF
RRRRCRRMH8RVR;
RRRRRR--l0kDH$bD
RRRRsRRVOsN0=R:RNVsOR0D*sRVNsO0;RRRRRRRRR--v0kDH$bDRC0ERNVsOF0HMR
RRRRR-N-R808RECCRGMbFC#M0
RRRRsRRCFGbM=R:R#sCHRxC5bCGF,MDRGsCb'FMDoCM0RE2+GRCbsFMR#-RE0HV$RR+4R;
RRRRRH#EVR0G:s=RCFGbMRR-CFGbM
O;RRRRRVRHRH#EVR0G<VR-s0NODH'Eo0ERE
CMRRRRRRRRsbCGFRM.:s=RCx#HCCR5GMbFOs,RCFGbMD.'C0MoE
2;RRRRRRRRVOsN0ROR:"=Rj&"RRNVsO;0G
RRRRRRRRNVsOR0#RR:=5EF0CRs#='>Rj;'2
RRRRRRRRH#0OR	$RR:=F5sRsNVsO;02
RRRRCRRDV#HRH#EVR0G<RRj0MEC
RRRRRRRRH#EVR0G:-=RRH#EV;0G
RRRRRRRRNVsOR0#:#=RE0HV_osHE50RsNVsO50RsNVsOE0'HRoE8MFI0sFRVOsN0H'EoRE
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-VOsN0D#'C0MoE2+4,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR_0FHCM0o5Cs#VEH02G2;R
RRRRRRsRVNOO0RRRR:"=Rj&"RRNVsO;0G
RRRRRRRRGsCb.FMR:RR=CRs#CHxRG5CbOFM,CRsGMbF.C'DMEo02R;
RRRRRDRRCsV0H0oERR:=V#NDCR;
RRRRR
RRRRRRRRRR-C-)I0sHCER0CFRVDIDFHRMo0RIFDCHM#VRFR8OFCFR0R	lNC$R#MC0E#NHxLRDC5FNPHC8RsssFR$#NH
MoRRRRRRRR-M-RFOM-F0M#NRM0HCM8GMRHRH#DOLCRCkON#FCRV#R"E0HVGR"RReRhZ-R4m-O0jRg
RRRRR-RR-H#0OR	$:F=RssR5VOsN00R5FM_H0CCosE5#HGV02V+ss0NO'oEHER
RRRRRR-R-RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RRRNVsO'0#DoCM08ERF0IMF2Rj2R;
RRRRR#RR00NsHR8G:0=RFM_H0CCosE5#HGV02V+ss0NO'oEHERR-VOsN0D#'C0MoER;
RRRRR#RR0	HO$=R:R''j;R
RRRRRRFRVsRRQHsMRVOsN0Q']t8]RF0IMFRRjDbFF
RRRRRRRRRRRRRHVQ=R<RN#0s80HGER0CRM
RRRRRRRRRRRRR#RR0	HO$=R:RH#0OR	$FssRVOsN025Q;R
RRRRRRRRRRMRC8VRH;RR
RRRRRCRRMD8RF;Fb
RRRRRRRRR--CRM8FsVRCHIs0RC
RRRRR#CDH#VRE0HVGRR=jER0CRM
RRRRRsRRCFGbM:.R=CRs#CHxRG5CbOFM,CRsGMbF.C'DMEo02R;
RRRRR#RR0	HO$:RR=sRFRV5ss0NORV5ss0NO'oEHERR-VOsN0DO'C0MoEFR8IFM0R2j2;R
RRRRRRVRHRssVNRO05ssVN'O0EEHoRI8FMR0FsNVsOE0'HRoE-sRVNOO0'MDCo+0E4>2RRNVsO
0GRRRRRRRR0MEC
RRRRRRRRVRRs0NOO=R:R""jRV&Rs0NOGR;
RRRRRRRRRNVsOR0#:s=RVOsN0sR5VOsN0H'Eo8ERF0IMFVRss0NO'oEHER
RRRRRRRRRRRRRRRRRRRRRRRRRRRR-VOsN0D#'C0MoE2+4;R
RRRRRRRRRD0CVsEHo0=R:RDVN#
C;RRRRRRRRCCD#
RRRRRRRRVRRs0NOO=R:RssVNRO05ssVN'O0EEHoRI8FMR0FsNVsOE0'H
oERRRRRRRRRRRRRRRRRRRRRRRRRRRR-sRVNOO0'MDCo+0E4
2;RRRRRRRRRsRVN#O0RRRR:"=Rj&"RRNVsO;0G
RRRRRRRRDRRCsV0H0oERR:=0Csk;R
RRRRRRMRC8VRH;R
RRRRRCHD#VER#HGV0RV>Rs0NOGH'Eo0ERE
CMRRRRRRRRsbCGFRM.R=R:RGsCb;FM
RRRRRRRRNVsOR0#R:RR=FR50sEC#>R=R''j2R;
RRRRRVRRs0NOORRRRR:=sNVsO50RsNVsOE0'HRoE8MFI0sFRVOsN0H'Eo-ERRNVsO'0ODoCM04E+2R;
RRRRRDRRCsV0H0oERR:=0Csk;R
RRRRRR0R#H$O	RR:=F5sRVOsN0&GRRssVNRO05ssVN'O0EEHoRV-Rs0NOOC'DMEo0
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRF0IMF2Rj2R;
RRRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-sRVNGO0'oEHERR>#VEH0>GRRRj
RRRRRsRRCFGbMR.RRR:=sbCGF
M;RRRRRRRRVOsN0R#RR=R:R""jR#&RE0HV_osHE50RVOsN0RG,0HF_Mo0CC5sR#VEH02G2;R
RRRRRRsRVNOO0RRRR:s=RVOsN0sR5VOsN0H'Eo8ERF0IMFVRss0NO'oEHERR-VOsN0DO'C0MoE2+4;R
RRRRRRCRDVH0soRE0:0=Rs;kC
RRRRRRRRR
RRRRRR-R-)sCIHR0C0RECVDFDFMIHoIR0FHRDMRC#FOVRFR8C0lFRNR	C#0$MEHC#xDNLCNR5P8FHRsCsF#sRNM$HoR
RRRRRR-R-RMMF-MOF#M0N0MRH8RCGH#MRDCHOROLCNCk#RRFV"H#EV"0GRRRRhReZ4O-m0g-j
RRRRRRRR#--0	HO$=R:RRFs5NVsOR0G5_0FHCM0oRCs5H#EV20GRI8FMR0FjR2
RRRRR-RR-RRRRRRRRRRRRRRRRRRRR&RRRssVNRO05ssVN'O0EEHoRV-Rs0NOOC'DMEo0RI8FMR0Fj;22
RRRRRRRRN#0s80HG=R:R_0FHCM0oRCs5H#EV20G;R
RRRRRR0R#H$O	RR:=';j'
RRRRRRRRsVFRHQRMsRVNGO0't]Q]FR8IFM0RDjRF
FbRRRRRRRRRRRRHQVRRR<=#s0N0GH8RC0EMR
RRRRRRRRRRRRRR0R#H$O	RR:=#O0H	F$RssRVNGO05;Q2
RRRRRRRRRRRR8CMR;HVRR
RRRRRRMRC8FRDF
b;RRRRRRRR
RRRRRRRRR--hRFI80FREsCRH0oERMEN8HR#8FCRVER0CsRFHMoHNODRFNMO0GRCb#sC#MHFReRhZ-R4m-O0jRg
RRRRR#RR0	HO$=R:RH#0OR	$F5sRF5sRsNVsO50RsNVsOE0'HRoE-sRVNOO0'MDCoR0E8MFI0jFR2;22
RRRRRRRRR--CRM8FsVRCHIs0RC
RRRRR8CMR;HV
RRRRVRRs0NO#jR52=R:RNVsOR0#5Rj2F#sR0	HO$R;R-m-RsER0C0R#H$O	R0LHR0HMFER0C1RpAR
RRRRRHVVRbH_#o=MRR_0FX5j4O'5OEEHo202RE
CMRRRRRRRRkNVsOR0R:V=Rs0NOORR+VOsN0
#;RRRRRRRRV#b_HRoM:V=RbH_#o
M;RRRRRDRC#RCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-#-RH#oMRCNsRV8HVCCsMR0
RRRRRkRRVOsN0=R:RNVsOR0O-sRVN#O0;RRRR-RR-DRNI#N$R#bFHP0HCCRs#0kD
RRRRRRRRRHVD0CVsEHo0ER0CRMRRRRRRRRRRRRRRR--wkHosFCRkI0REEHORo#HMFR0RCk#
RRRRRRRRVRRbH_#o:MR=bRV_o#HMR;
RRRRRCRRD
#CRRRRRRRRRbRV_o#HM=R:ROO5'oEHE
2;RRRRRRRRCRM8H
V;RRRRRMRC8VRH;R
RRRRR-M-RFNslDCHx
RRRRVRRb#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>kNVsO
0,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=s>RCFGbM
.,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRo#HMRRRRRRRRRRR=V>RbH_#o
M,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRH#0OR	$RRRRRRRR=#>R0	HO$R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRoRMk8NsRRRRRRRRRR=>oskN8
2;RRRRCRM8H
V;RRRRskC0sVMRb#sCk;D0
CRRMV8Rk0MOHRFMl;NO
R
R-"-Rs"ClRMVkOF0HMR
RVOkM0MHFRlsCN8HMC5sR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRRRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRNoksR8RRRRRRh:Rq)azqRpRR=R:RFVDNo0_k8Ns_0LH#R;R-M-RkClLsVRFRNoksL8RH
0#RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs;RR--OOEC	FRVssRCs#Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0RERRh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0ERRR:hzqa)Rqp:l=RNlGHkDl5'oEHEs,R'oEHER2;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRMOF#M0N0HR8PNoksR8RRRRRR:RRRahqzp)qRR:=oskN8R;R-8-RH#PHHRFMoskN8HRL0R#
RPRRNNsHLRDCD0Vb$,bCRbsV0C$bRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDVCRb#sCkRD0RRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RRRRPHNsNCLDRVkDs0NO,sRkVOsN0RR:zQh1t7h Rs5VNHO0FIM_HE80RI8FMR0Fj
2;RRRRPHNsNCLDRNVsO,0sRNVsOR0DRRR:zQh1t7h Rs5VNHO0FIM_HE80+P8HoskN8FR8IFM0R;j2R-R-RosHER0
RPRRNNsHLRDCsNVsOR0RRRRRRRRRRz:Rht1QhR 75NVsO'0ssoNMCR2;R-RR-CRs#0kDRNVsOF0HMR
RRNRPsLHND#CRVOsN0RRRRRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH08E+HkPoNRs88MFI0jFR2R;R-s-RCD#k0sRVNHO0FRM
RPRRNNsHLRDCCFGbMRD,CFGbMRsRR1:RQ th7CR5GMbFC_M0I0H8ER-48MFI0jFR2R;R-C-RGMbFC#M0
RRRRsPNHDNLCCRsGMbFRRRRRRRRR:RRRt1QhR 75bCGFMMC0H_I8R0E8MFI0jFR2R;R-s-RCD#k0GRCbCFMMR0
RPRRNNsHLRDCV#b_HRoMRRRRRRRRR1:Raz7_pQmtBR;RRRRRR-R-Ro#HMVRFR#sCk
D0RRRRPHNsNCLDRH#EVR0$RRRRRRRRRRR:Q hat; )RRRRRRRRR-RR-CR8MlFsNMDRkClLsER#H
V0RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RLHCoM-RR-CRslMNH8
CsRRRRH5VRVOsN0MHF_8IH0=ERRFjRs'RDDoCM0<ERRF(Rs'RsDoCM0<ERRR(20MEC
RRRRDRRV$b0b:CR=#RHGR;
RCRRD
#CRRRRRVRDbb0$C=R:RNOD#b#VR,5DRCOEOC	_sssF2R;
RRRRRbsV0C$bRR:=O#DN#RVb5Rs,OOEC	s_Cs2Fs;R
RRMRC8VRH;R
RRVRHRV5Dbb0$CRR=HR#GFssRV$b0b=CRRGH#2ER0CRM
RRRRRsVbCD#k0=R:R05FE#CsRR=>'2X';R
RRDRC#RHV5bDV0C$bRM=RNFMRsVRDbb0$CRR=JCkH0N_MMR2
RRRRRRFs5bsV0C$bRM=RNFMRsVRsbb0$CRR=JCkH0N_MMR2
RRRRRR--)kC0sJMRk0HCRhhq, RQ 6 (cg-4U(6-344,
RRRRFRRsDR5V$b0b=CRR#bF_VHMRRFsD0Vb$RbC=CRMoM_HVR2R-H-RMsVRCGlR
RRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,R6
RRRRRRFs5bsV0C$bRb=RFx#_CRsFFssRV$b0b=CRRoMC_sxCF02RERCMR-RR-RRGsRCljR
RRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,6RRRRRbRVskC#D:0R=MRJNbMVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRR#CDH5VRs0Vb$RbC=FRb#M_HVsRFRbsV0C$bRM=RCHo_MRV20MECRRRRRR--GCRslMRHVRR=jR
RRRRRVCbs#0kDRR:=xFCsV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RCRRDV#HRL5N#25DRN<RLs#5202RE
CMRRRRRbRVskC#D:0R=;RD
RRRR#CDCR
RRRRRV#b_HRoM:0=RFj_X455DDH'Eo2E2;RRRR-R-Ro#HMR
RRRRRD#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4D
2,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRRbDV0C$bRR:=O#DN#RVb5CDs#CHx,NRVD2#C;RRRRRRRR-R-RsCsFRs#NCDsNR8$OOEC	
C8RRRRRsRsCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425s,R
RRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRsRRV$b0b:CR=DRONV##bsR5sHC#xRC,V#NDCR2;RRRRRRRR-C-RsssF#DRNs8CN$EROCCO	8R
RRRRRVOsN0RDR:5=RFC0Es=#R>jR''
2;RRRRRsRLC_N	MLklC5sR
RRRRRRRRoNsRRRRRRRRRR=>D#sCH,xC
RRRRRRRR0Vb$RbRRRRRRR=>D0Vb$,bC
RRRRRRRRM8CFNslDCHxRR=>8FCMsDlNH,xC
RRRRRRRRNVsOR0RRRRRRR=>ksDVN,O0
RRRRRRRRbCGFRMRRRRRRR=>CFGbM;D2
RRRRVRRs0NODVR5s0NOH_FMI0H8EH+8PNoks88RF0IMFHR8PNoksR82:k=RDNVsO
0;RRRRR-R-RosHE#0RH
8CRRRRRsRVNsO0RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR:RR=FR50sEC#>R=R''j2R;
RRRRRCLsNM	_kClLs
R5RRRRRRRRNRsoRRRRRRRR=s>RsHC#x
C,RRRRRRRRV$b0bRRRRRRR=s>RV$b0b
C,RRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx
C,RRRRRRRRVOsN0RRRRRRR=k>RsNVsO
0,RRRRRRRRCFGbMRRRRRRR=C>RGMbFs
2;RRRRRsRVNsO0Rs5VNHO0FIM_HE80+P8HoskN8FR8IFM0RP8HoskN8:2R=sRkVOsN0R;
RRRRRGsCbRFMRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=R:RG5CbsFM5bCGF'MsEEHo2G&CbsFM2R;
RRRRRH#EVR0$RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR=R:R_0FHCM0o5CsCFGbM-DRRGsCb2FM;R
RRRRRH5VR#VEH0>$RRRj20MEC
RRRRRRRRNVsOR0s:#=RE0HV_osHE50RVOsN0Rs,#VEH0;$2
RRRRRRRRGsCbRFM:s=RCFGbMRR+#VEH0
$;RRRRRMRC8VRH;R
RRRRRH5VRVOsN0/sR=2RjRC0EMR
RRRRRR-R-RlsC
RRRRRRRRssVNRO0:V=Rs0NODCRslsRVNsO0;RRRRR--kHM#o8MCRlsC
RRRRRRRRs#VNRO0:s=RVOsN0#R5VOsN0N'sM2oC;RRRRRRRRRRR-D-RFsICR0LH#R
RRRRRR-R-RsMFlHNDxRC
RRRRRVRRb#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>#NVsO
0,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFRRRRRRRRR>R=RGsCb,FM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR#MHoRRRRRRRRR=RR>bRV_o#HMR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRMNoksR8RRRRRR=RR>HR8PNoks;82
RRRRCRRD
#CRRRRRRRR-Q-RVCRIRH#EV"0RVOsN0Rs"#VFRN0sRERN0HL0RClOFCx#RC,sFR0sCkRsMxFCs3R
RRRRRRbRVskC#D:0R=CRxsbFVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRR8CMR;HV
RRRR8CMR;HV
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFRlsCN8HMC
s;
-RR-lR"FR8"VOkM0MHF
VRRk0MOHRFMlkF8D5FR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0oskN8RRRRRRR:qRhaqz)pRRRRR:=VNDF0k_oN_s8L#H0;-RR-kRMlsLCRRFVoskN8HRL0R#
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRFROMN#0MV0Rs0NOH_FMI0H8ERRR:qRhaqz)p=R:Rl-RH5MCDF'DIs,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0ERRR:hzqa)Rqp:l=RNlGHkDl5'oEHEs,R'oEHER2;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRsPNHDNLCVRDbb0$Cs,RV$b0b:CRRDPNHV8_bN#00
C;RRRRPHNsNCLDRsVbCD#k0RRRRRRRRRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RRNRPsLHNDsCRCCls#RRRRRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RCRLoRHMRR--sNClHCM8sR
RRVRHRs5VNHO0FIM_HE80Rj=RRRFsDC'DMEo0R(<RRRFssC'DMEo0R(<R2ER0CRM
RRRRRbDV0C$bRR:=H;#G
RRRR#CDCR
RRRRRD0Vb$RbC:O=RD#N#V5bRDO,RE	CO_sCsF;s2
RRRRsRRV$b0b:CR=DRONV##bsR5,EROC_O	CFsss
2;RRRRCRM8H
V;RRRRH5VRD0Vb$RbC=#RHGsRFRbsV0C$bRH=R#RG20MEC
RRRRVRRb#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRCHD#VDR5V$b0b=CRRMMNRRFsD0Vb$RbC=kRJH_C0M2NM
RRRRFRRssR5V$b0b=CRRMMNRRFss0Vb$RbC=kRJH_C0M2NM
RRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,R4
RRRRRRFs5bDV0C$bRb=RFH#_MFVRsVRDbb0$CRR=M_CoH2MVRRRRRRRRR-RR-MRHVCRsl
RGRRRRR-R-R0)CkRsMJCkH0qRhhQ,R (  64c-g-U6(,346R
RRRRRF5sRs0Vb$RbC=FRb#C_xsFFRsVRsbb0$CRR=M_CoxFCs2ER0CRMRR-R-RsGRCjlR
RRRR-RR-CR)0MksRHJkCh0RqRh,Q   (-6c46gU-4(3,R6
RRRRRsVbCD#k0=R:RNJMMRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRCHD#VsR5V$b0b=CRR#bF_VHMRRFss0Vb$RbC=CRMoM_HV02RERCMRRRR-G-RRlsCRVHMRj=R
RRRRVRRb#sCkRD0:x=RCVsFbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I820E;R
RRDRC#RC
RRRRRlsCsRC#:s=RCHlNMs8CRR5DRRRRRRRRR>R=R#NL5,D2
RRRRRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=N>RLs#52R,
RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$C>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRNoksR8RRRRRRR=>oskN8R,
RRRRRRRRRRRRRRRRRRRRRRRRREROC_O	CFsss>R=RDVN#
C,RRRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDx=CR>CR8MlFsNxDHC
2;RRRRR-R-R7vmRRH#0REC#CNlRRN#), vR0LkRk$FRR8F#CFl0MEHoHR8VsVCCRM0IEH0
RRRR-RR-CRMoHN0PPCRNCDk#R
RRRRRH5VRHM#_C0oNHRPC52D2RC0EMR
RRRRRRCRsl#sCRR:=-CRsl#sC;R
RRRRRCRM8H
V;RRRRRVRHR#5H_oMCNP0HCDR52RR=HM#_C0oNHRPC5Rs2FssRCCls#RR=j02RE
CMRRRRRRRRVCbs#0kDRR:=ssClC
#;RRRRRDRC#RC
RRRRRVRRb#sCkRD0:N=R858RDRRRRRRRRRRR=s>RCCls#R,
RRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=s>R,R
RRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRoskN8RRRRRRR=o>Rk8Ns,R
RRRRRRRRRRRRRRRRRRRRRRORRE	CO_sCsF=sR>NRVD,#C
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx2R;RRRRRRRR
RRRRR8CMR;HV
RRRR8CMR;HV
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFR8lFk;DF
R
R-1-RJskNCFRsFF0RVRRNVNDF0oHMRHbFMM0RkClLsR3R7CFMRHk#MhoRCFI0MR'#Qs0CNF0HMR3
RMVkOF0HMJR#s50R
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRRRRRRRR--VNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DC
RRRRMOF#M0N0kRoNRs8RRRRRRR:hzqa)RqpR:RR=DRVF_N0oskN8H_L0
#;RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDx
C2RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=kRoN-s8N'soD;FIR-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)Rqp:N=RsEo'H;oER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHND#CRHRoMRRRRRRRRRRR:1_a7ztpmQ
B;RRRRPHNsNCLDRsVbCD#k0RRRRRRR:DRVFRN05oNs'MsNo;C2
RRRRsPNHDNLCbRV0C$bRRRRRRRRRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDHCRCFGbMRRRRRRRRRR:1hQt C75GMbFC_M0I0H8ER-48MFI0jFR2R;R-C-RGMbFC#M0
RRRRsPNHDNLCGRCbRFMRRRRRRRRR1:RQ th7G5CbCFMMI0_HE80RI8FMR0FjR2;R-RR-GRCbCFMM
0#RRRRPHNsNCLDRNkVOR0RRRRRRRRR:VRkH8GCRR5j8MFI0NFRsDo'F;I2
RRRRsPNHDNLCNRVOR0RRRRRRRRRRk:RVCHG8.R5RI8FMR0F-NVsOF0HMH_I820E;-RR-sRVNHO0FRM
RPRRNNsHLRDCsLC#RRRRRRRRR:RRRHkVGRC85OVN0H'Eo4E+RI8FMR0FV0NO'IDF2R;
RoLCHRMR-#-RJskNCFRsFR0
RVRRbb0$C=R:RNBD#b#VRs5NoO,RE	CO_sCsF;s2
RRRRNOD#N#O#:CRR#ONCbRV0C$bR
H#RRRRRERICHMR#=GR>R
RRRRRRbRVskC#D:0R=FR50sEC#>R=R''X2R;
RRRRRCIEMNRMMRR|JCkH0N_MM
R|RRRRRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,4RRRRRRRRM_CoMlFsN|DRRoMC_M8CFNslDRR|M_CoHRMV=R>RRRRR-#-RJRs05oMC2R
RRRRRR-R-R0)CkRsMJCkH0qRhhQ,R (  64c-g-U6(334nR
RRRRRRbRVskC#D:0R=MRJNbMVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0oE-k8Ns,R
RRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRIRRERCMb_F#HRMV=R>RRRRRRRRRRRRRRRRRRR--10JsRM5HVR2,skC0sHMRMMVHH
0$RRRRRRRRVCbs#0kDRR:=b_F#HVMVbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8-0EoskN8R,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRIRRERCMb_F#xFCsRR=>RRRRRRRRRRRRRRRRRR--skC0sjMR
RRRRRRRRsVbCD#k0=R:RsxCFRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8Ek-oN,s8
RRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRERICMMRCxo_CRsF=R>RRRRRRRRRRRRRRRRR-Q-R (  64c-g-U6nR3dskC0s-MRjR
RRRRRRbRVskC#D:0R=CRMoC_xsbFVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0oE-k8Ns,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRIRRERCMFC0Es=#R>R
RRRRRRsRLC_N	MLklC5sRNRsoRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRROOEC	s_CsRFs=V>RNCD#,R
RRRRRRRRRRRRRRRRRRRRRVOsN0RRRRRRR=k>RV0NO,R
RRRRRRRRRRRRRRRRRRRRRCFGbMRRRRRRR=H>RCFGbMR,
RRRRRRRRRRRRRRRRRRRRRo#HMRRRRRRRRR=>#MHo2R;
RRRRRCRRGMbFRR:=sHC#x5CRHbCGF4M+,GRCb'FMDoCM0;E2R-RR-CRo0GRCbCFMMR0
RRRRRVRRNRO0RR:=sHC#x5CRkOVN0V,RN'O0EEHo,NRVOD0'F;I2
RRRRRRRRRHV5bCGFjM52RR='24'RC0EMR
RRRRRRRRRV0NORR:=V0NORN#DRR4;RRRRRRRRR-R-R.*R3Rj
RRRRRCRRMH8RVR;
RRRRRCRRGMbFRR:=#VEH0H_soRE05bCGFRM,4R2;RRRRRRRRR-RR-GRCbCFMM.0/
RRRRRRRRR--h0CIF#M'RCH0sHN0F-MRRFsF0=R:RR54+sRNo/2RRR.
RRRRRsRRCR#LRR:=5OVN0RR+4#2Rs4NR;R
RRRRRRFRVsRR[HjMRRR0FVOsN0MHF_8IH0cE/RFDFbR
RRRRRRRRR-R-RRFsF0=R:RF5sF+0RRs5NoF/sF202/R.
RRRRRRRRR#sCL=R:R#sCHRxC5oNsRRRRRRRRRRRR=5>RsLC#R5+RV0NO/#sCLR22#RsN4R,
RRRRRRRRRRRRRRRRRRRRRRRRRVDC0M_H8RCGRRRR=s>RC'#LEEHo,R
RRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>CRs#DL'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>VCHG8s_0kNMO0
C,RRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>VCHG8s_IN;b2
RRRRRRRR8CMRFDFbR;
RRRRRVRRb#sCkRD0:M=RFNslDCHxRs5VNRO0RRRRRRRRRR=>sLC#,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFRMRRRRRRRRR=C>RGMbF-
4,RRRRRRRRRRRRRRRRRRRRRRRRRRRRR#RRHRoMRRRRRRRRR>R=R''j,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=N>RsEo'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>NR-sDo'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRMRRoskN8RRRRRRRR>R=RNoks;82
RRRR8CMR#ONCDRONO##N;#C
RRRR0sCkRsMVCbs#0kD;R
RCRM8VOkM0MHFRs#J0
;
RkRVMHO0FQMR#C_hoHN0P5CRNRso:hRz)m 1p7e _FVDNR02skC0sAMRm mpqHhR#R
RR-R-ROaCEOMHN$DDRR-j#kEFDs8RCs0kMVR"NCD#"L,RkQ0R'DlRCHNPM0oRERN0OCN#R0Fk3R
RLHCoMR
RRCRs0MksRF50_4Gj5oNs5oNs'oEHER22=4R''
2;RMRC8kRVMHO0FQMR#C_hoHN0P
C;
-RR-FROlsbNCkRVMHO0F
M#R-R-RR=,/R=,>R=,<R=,<>,R
R
RVOkM0MHFRRCJ5RRRRRRRRRRRRRRRRRRRRRRRR-R-RkCJN=DR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpq:hR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMApmm 
qhR#RH
RRRRsPNHDNLCVRDbb0$Cs,RV$b0bRCRRRRRRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDHCR#J_Ck,NDR_H#ksMF8CCs8RR:Apmm ;qh
RRRRMOF#M0N0sRVNHO0FIM_HE80RRRRRRRRRh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0ERRRRRRRR:qRhaqz)p=R:RGlNHllk5ED'H,oEREs'H2oE;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RPRRNNsHLRDCD#sCH,xCRCss#CHxRRRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RoLCHRMR-C-RJDkN
RRRRRHV5NVsOF0HMH_I8R0E=RRjFDsR'MDCoR0E<RR(FssR'MDCoR0E<2R(RC0EMR
RRRRRskC0sVMRNCD#;R
RRDRC#RC
RRRRRbDV0C$bRR:=O#DN#RVb5RD,OOEC	s_Cs2Fs;R
RRRRRs0Vb$RbC:O=RD#N#V5bRsO,RE	CO_sCsF;s2
RRRR8CMR;HV
RRRRRHV5bDV0C$bRM=RCxo_CRsFFDsRV$b0b=CRR#bF_sxCFN2RMR8
RRRRRV5sbb0$CRR=M_CoxFCsRRFss0Vb$RbC=FRb#C_xsRF20MEC
RRRRHRR#J_CkRND:0=Rs;kC
RRRR#CDCR
RRRRRD#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4D
2,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRRCss#CHxRR:=sHC#x5CRNRsoRRRRRRRRR=RR>FR0_4Gj5,s2
RRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNH_xCH=MR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHC
2;RRRRR#RH_kCJN:DR=0R5FD_#Ps5DCx#HC=2RR_0F#5DPs#sCH2xC2R;
RCRRMH8RVR;
RHRRVOR5E	CO_sCsFRs20MEC
RRRRHRR#M_kFCs8sRC8:z=RM8FsC8sCRR5G=D>R,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$RRRR=>s
2;RRRRCCD#
RRRRHRR#M_kFCs8sRC8:V=RNCD#;R
RRMRC8VRH;R
RRCRs0MksR_H#CNJkDMRN8FRM0#RH_FkMss8CC
8;RMRC8kRVMHO0FCMRJ
;
RkRVMHO0FDMR0RR5RRRRRRRRRRRRRRRRRRRRRRRR-D-RCR##0MENRR<
RDRR,RRsRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RRRRRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpq:hR=DRVF_N0OOEC	s_Cs;Fs
RRRRMOF#M0N0CR8MlFsNxDHCRR:Apmm Rqh:V=RD0FN_M8CFNslDCHx2R
RRCRs0MksRmAmph q
HRR#R
RRFROMN#0MV0Rs0NOH_FMI0H8ERRRRRRRRRRRRRR:hzqa)Rqp:-=RlCHM5DD'FRI,sF'DIR2;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0GRCbCFMMI0_HE80RRRRRRRRRRRRRh:Rq)azq:pR=NRlGkHll'5DEEHo,'RsEEHo2R;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRPHNsNCLDRbDV0C$b,VRsbb0$CRRRRRRRRRRR:NRPD_H8V0b#N;0C
RRRRsPNHDNLCGRCbRD,CsGbRRRRRRRRRRRRRRRRRz:Rht1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2
RRRRsPNHDNLCsRVNDO0,sRVNsO0RRRRRRRRRRRRRz:Rht1QhR 75NVsOF0HMH_I8-0E4FR8IFM0R;j2
RRRRsPNHDNLC#RH_#DC#E_0NRM,Hk#_M8FsC8sCRA:Rm mpq
h;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRRRRRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RCRLo
HMRRRRH5VRVOsN0MHF_8IH0=ERRFjRs'RDDoCM0<ERRF(Rs'RsDoCM0<ERRR(20MEC
RRRRHRR#C_D#0#_ERNM:V=RNCD#;R
RRDRC#RC
RRRRRCDs#CHxRR:=sHC#x5CRNRsoRRRRRRRRR=RR>FR0_4Gj5,D2
RRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNH_xCH=MR>CR8MlFsNxDHCR,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHC
2;RRRRRsRsCx#HC=R:R#sCHRxC5oNsRRRRRRRRRRRR=0>RFj_G425s,R
RRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRHRRVFR0_4Gj5DD5'oEHER22=FR0_4Gj5ss5'oEHER220MECR-R-Ro#HMHRL0R#
RRRRRCRRGRbD:z=Rht1Qh5 7D#sCH5xCCFGbM0CM_8IH04E-RI8FMR0Fj;22
RRRRRRRRbCGs=R:R1zhQ th7s5sCx#HCG5CbCFMMI0_HE80-84RF0IMF2Rj2R;
RRRRRHRRVGRCb=DRRbCGsER0CRM
RRRRRRRRRNVsOR0D:z=Rht1QhR 75_0F#5DPD#sCH5xC-84RF0IMFVR-s0NOH_FMI0H8E222;R
RRRRRRRRRVOsN0:sR=hRz1hQt 57R0#F_DsP5sHC#x-C54FR8IFM0Rs-VNHO0FIM_HE802;22
RRRRRRRRHRRVFR0_4Gj5DD5'oEHER22=jR''ER0CRMRRRRRRRRRR-R-R#bFHP0HCkRMlsLC
RRRRRRRRRRRR_H#D#C#_N0EM=R:Rs5VNDO0RV<Rs0NOs
2;RRRRRRRRRDRC#RC
RRRRRRRRRHRR#C_D#0#_ERNM:5=RVOsN0>DRRNVsO20s;RRRRRRR-M-RC0oNH
PCRRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRRRHV0GF_jD455ED'H2oE2RR='Rj'0MECRRRRRRRRRRRR-b-RF0#HHRPCMLklCRs
RRRRRRRRRHRR#C_D#0#_ERNM:5=RCDGbRC<RG2bs;R
RRRRRRRRRCCD#
RRRRRRRRRRRR_H#D#C#_N0EM=R:RG5Cb>DRRbCGsR2;RRRRRRRRR-R-RoMCNP0HCR
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8H
V;RRRRRDRC#RC
RRRRRDRRV$b0b:CR=DRONV##bDR5,EROC_O	CFsss
2;RRRRRRRRs0Vb$RbC:O=RD#N#V5bRsO,RE	CO_sCsF;s2
RRRRRRRRRHV5bDV0C$bRM=RCxo_CRsFNRM8s0Vb$RbC=FRb#C_xsRF20MEC
RRRRRRRRHRR#C_D#0#_ERNM:V=RNCD#;RRRRRRRRR---<jRRsjRCs0kMV#RNCD#3R
RRRRRRDRC#RC
RRRRRRRRR_H#D#C#_N0EM=R:RF50_4Gj5DD5'oEHER22>FR0_4Gj5ss5'oEHE222;R
RRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RRRRHOVRE	CO_sCsF0sRE
CMRRRRR#RH_FkMss8CC:8R=MRzFCs8sRC85=GR>,RD
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$=s>R2R;
RCRRD
#CRRRRR#RH_FkMss8CC:8R=NRVD;#C
RRRR8CMR;HV
RRRR0sCkRsMHD#_C_##0MENR8NMR0MFR_H#ksMF8CCs8R;
R8CMRMVkOF0HM0RD;R

RMVkOF0HM0RoRR5RRRRRRRRRRRRRRRRRRRRRR-RR-sRoCCN0sER0N>MR
RRRRRD,sRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp h=R:RFVDNO0_E	CO_sCsF
s;RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpq:hR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMApmm 
qhR#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80R:RRRahqzp)qRR:=-MlHC'5DD,FIRDs'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERRR:qRhaqz)p=R:RGlNHllk5ED'H,oEREs'H2oE;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RPRRNNsHLRDCD0Vb$,bCRbsV0C$bRP:RN8DH_#Vb0CN0;R
RRNRPsLHNDCCRG,bDRbCGsRRRRRRR:hRz1hQt 57RCFGbM0CM_8IH04E-RI8FMR0Fj
2;RRRRPHNsNCLDRNVsO,0DRNVsOR0sRRR:zQh1t7h Rs5VNHO0FIM_HE80-84RF0IMF2Rj;R
RRNRPsLHNDHCR#s_oCCN0sE_0NRMR:mRAmqp hR;
RPRRNNsHLRDCHk#_M8FsC8sCRRRRRA:Rm mpq
h;RRRRPHNsNCLDRCDs#CHx,sRsCx#HCRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RLHCoM-RR-sRoCCN0sE_0NRM
RHRRVVR5s0NOH_FMI0H8ERR=jsRFRDD'C0MoERR<(sRFRDs'C0MoERR<(02RE
CMRRRRR#RH_CosNs0C_N0EM=R:RDVN#
C;RRRRCCD#
RRRRDRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>0GF_jD452R,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRs#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R_0FG5j4s
2,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRRRHV0GF_jD455ED'H2oE2RR=0GF_js455Es'H2oE2ER0CRMRRRRRRRRRRRRR-#-RHRoML#H0
RRRRRRRRbCGD=R:R1zhQ th7s5DCx#HCG5CbCFMMI0_HE80-84RF0IMF2Rj2R;
RRRRRCRRGRbs:z=Rht1Qh5 7s#sCH5xCCFGbM0CM_8IH04E-RI8FMR0Fj;22
RRRRRRRRRHVCDGbRC=RGRbs0MEC
RRRRRRRRVRRs0NOD=R:R1zhQ th70R5FD_#Ps5DCx#HC45-RI8FMR0F-NVsOF0HMH_I820E2
2;RRRRRRRRRsRVNsO0RR:=zQh1t7h RF50_P#D5Css#CHx5R-48MFI0-FRVOsN0MHF_8IH02E22R;
RRRRRRRRRRHV0GF_jD455ED'H2oE2RR='Rj'0MECRRRRRR--bHF#0CHPRlMkL
CsRRRRRRRRRRRRHo#_s0CNC0s_ERNM:V=Rs0NODRR>VOsN0
s;RRRRRRRRRDRC#RC
RRRRRRRRRHRR#s_oCCN0sE_0N:MR=sRVNDO0RV<Rs0NOsR;RRRRRRRRRRRRRRRRR-M-RC0oNH
PCRRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRRRHV0GF_jD455ED'H2oE2RR='Rj'0MECRRRRRR--bHF#0CHPRlMkL
CsRRRRRRRRRRRRHo#_s0CNC0s_ERNM:C=RGRbD>GRCb
s;RRRRRRRRRDRC#RC
RRRRRRRRRHRR#s_oCCN0sE_0N:MR=GRCb<DRRbCGsR;RRR--MNCo0CHP
RRRRRRRRCRRMH8RVR;
RRRRRCRRMH8RVR;
RRRRR#CDCR
RRRRRRVRDbb0$C=R:RNOD#b#VR,5DRCOEOC	_sssF2R;
RRRRRsRRV$b0b:CR=DRONV##bsR5,EROC_O	CFsss
2;RRRRRRRRH5VRD0Vb$RbC=FRb#C_xsNFRMs8RV$b0b=CRRoMC_sxCF02RE
CMRRRRRRRRR#RH_CosNs0C_N0EM=R:RDVN#RC;RRRR-j-RR->RjCRs0Mks#NRVD3#C
RRRRRRRR#CDCR
RRRRRRRRRHo#_s0CNC0s_ERNM:0=RFj_G455DDH'Eo2E2R0<RFj_G455ssH'Eo2E2;R
RRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRCRM8H
V;RRRRHOVRE	CO_sCsF0sRE
CMRRRRR#RH_FkMss8CC:8R=MRzFCs8sRC85=GR>,RD
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$=s>R2R;
RCRRD
#CRRRRR#RH_FkMss8CC:8R=NRVD;#C
RRRR8CMR;HV
RRRR0sCkRsMHo#_s0CNC0s_ERNMNRM8MRF0Hk#_M8FsC8sC;R
RCRM8VOkM0MHFR;o0
R
R-b-RkFsb#RC:/V=Rk0MOH
FMRkRVMHO0FMMRCRR5RRRRRRRRRRRRRRRRRRRRRRRR-M-RFC0RJDkNR
/=RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm Rqh:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMmRAmqp hR
RHR#
RPRRNNsHLRDCHC#_JDkN,#RH_FkMss8CC:8RRmAmph q;R
RLHCoMR
RR#RH_kCJN:DR=JRCRR5DRRRRRRRRR>R=R
D,RRRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=s>R,R
RRRRRRRRRRRRRRRRRREROC_O	CFsss>R=RDVN#
C,RRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx;C2
RRRRRHVOOEC	s_CsRFs0MEC
RRRRHRR#M_kFCs8sRC8:z=RM8FsC8sCRR5G=D>R,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$RRRR=>s
2;RRRRCCD#
RRRRHRR#M_kFCs8sRC8:V=RNCD#;R
RRMRC8VRH;R
RRCRs0MksR0MFR#5H_kCJNNDRMM8RFH0R#M_kFCs8s2C8;R
RCRM8VOkM0MHFR;MC
R
RVOkM0MHFRRDC5RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-D-RCR##0MENRRFsCNJkDFR0R
<=RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp h=R:RFVDN80_CsMFlHNDx
C2RRRRskC0sAMRm mpqRh
R
H#RRRRPHNsNCLDR_H#oNsC0_Cs0MEN,#RH_FkMss8CC:8RRmAmph q;R
RLHCoMR
RR#RH_CosNs0C_N0EM=R:RRo05RDRRRRRRRRRRR=>DR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRR>R=R
s,RRRRRRRRRRRRRRRRRRRRRRRRRORRE	CO_sCsF=sR>NRVD,#C
RRRRRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx;C2
RRRRRHVOOEC	s_CsRFs0MEC
RRRRHRR#M_kFCs8sRC8:z=RM8FsC8sCRR5G=D>R,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$RRRR=>s
2;RRRRCCD#
RRRRHRR#M_kFCs8sRC8:V=RNCD#;R
RRMRC8VRH;R
RRCRs0MksR0MFR_H#oNsC0_Cs0MENR8NMR0MFR_H#ksMF8CCs8R;
R8CMRMVkOF0HMCRD;R

RMVkOF0HMCRoRR5RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--oNsC0RCs0MENRRFsCNJkDFR0R
>=RRRRDs,RRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp h=R:RFVDN80_CsMFlHNDx
C2RRRRskC0sAMRm mpqRh
R
H#RRRRPHNsNCLDR_H#D#C#_N0EMH,R#M_kFCs8sRC8:mRAmqp hR;
RoLCHRM
RHRR#C_D#0#_ERNM:D=R0DR5RRRRRRRRR=RR>,RD
RRRRRRRRRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=>sR,
RRRRRRRRRRRRRRRRRRRRRORRE	CO_sCsF=sR>NRVD,#C
RRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRR=>8FCMsDlNH2xC;R
RRVRHRCOEOC	_sssFRC0EMR
RRRRRHk#_M8FsC8sCRR:=zsMF8CCs8GR5RR=>DR,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR$>R=R;s2
RRRR#CDCR
RRRRRHk#_M8FsC8sCRR:=V#NDCR;
RCRRMH8RVR;
RsRRCs0kMFRM0#RH_#DC#E_0NNMRMM8RFH0R#M_kFCs8s;C8
CRRMV8Rk0MOHRFMo
C;
VRRk0MOHRFM""?=R,5pR:)RR)zh p1me_ 7VNDF0s2RCs0kMaR17p_zmBtQR
H#RRRRO#FM00NMRNVsOF0HMH_I8R0ERRRRRRRR:qRhaqz)p=R:RH-lMDC5'IDF,'RsD2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0RERRRRRR:RRRahqzp)qRR:=lHNGl5klDH'EoRE,sH'Eo;E2R-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHNDDCRV$b0bRC,s0Vb$RbCRRRRRRR:PHND8b_V#00NCR;
RPRRNNsHLRDCHC#_JDkN,#RH_FkMss8CC:8RR71a_mzpt;QB
RRRRsPNHDNLCsRDCx#HCs,RsHC#xRCRRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
LRRCMoHR-R-R
?=RRRRH5VRVOsN0MHF_8IH0=ERRFjRs'RDDoCM0<ERRF(Rs'RsDoCM0<ERRR(20MEC
RRRRsRRCs0kMXR''R;
RCRRD
#CRRRRRVRDbb0$C=R:RNOD#b#VR,5DRFVDNO0_E	CO_sCsF;s2
RRRRsRRV$b0b:CR=DRONV##bsR5,DRVF_N0OOEC	s_Cs2Fs;R
RRMRC8VRH;R
RRVRHRV5Dbb0$CRR=M_CoxFCsRRFsD0Vb$RbC=FRb#C_xsRF2N
M8RRRRRsR5V$b0b=CRRoMC_sxCFsRFRbsV0C$bRb=RFx#_C2sFRC0EMR
RRRRRHC#_JDkNRR:=';4'
RRRR#CDCR
RRRRRD#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R
D,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RFVDN80_CsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=V>RD0FN_M8CFNslDCHx2R;
RRRRRCss#CHxRR:=sHC#x5CRNRsoRRRRRRRRR=RR>,Rs
RRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNH_xCH=MR>DRVF_N08FCMsDlNH,xC
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>VNDF0C_8MlFsNxDHC
2;RRRRR#RH_kCJN:DR=FR0_D#kPs5DCx#HC?2R=FR0_D#kPs5sCx#HC
2;RRRRCRM8H
V;RRRRH5VRVNDF0E_OC_O	CFsss02RE
CMRRRRRVRHRV5Dbb0$CRR=MRNMFDsRV$b0b=CRRHJkCM0_NFMRsR
RRRRRRRRRs0Vb$RbC=NRMMsRFRbsV0C$bRJ=Rk0HC_MMN2ER0CRM
RRRRRHRR#M_kFCs8sRC8:'=R4
';RRRRRDRC#RC
RRRRRHRR#M_kFCs8sRC8:'=Rj
';RRRRRMRC8VRH;R
RRDRC#RC
RRRRR_H#ksMF8CCs8=R:R''j;R
RRMRC8VRH;R
RRCRs0MksR_H#CNJkDMRN8FRM0#RH_FkMss8CC
8;RMRC8kRVMHO0F"MR?;="
R
RVOkM0MHFR/"?=5"Rp),RRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RRFROMN#0MV0Rs0NOH_FMI0H8ERRRRRRRRRR:hzqa)Rqp:-=RlCHM5DD'FRI,sF'DIR2;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0GRCbCFMMI0_HE80RRRRRRRRRh:Rq)azq:pR=NRlGkHll'5DEEHo,'RsEEHo2R;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRPHNsNCLDRbDV0C$b,VRsbb0$CRRRRRRR:NRPD_H8V0b#N;0C
RRRRsPNHDNLC#RH_kCJNRD,Hk#_M8FsC8sCR1:Raz7_pQmtBR;
RPRRNNsHLRDCD#sCH,xCRCss#CHxRRRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RoLCHRMR-?-R/R=
RHRRVVR5s0NOH_FMI0H8ERR=jsRFRDD'C0MoERR<(sRFRDs'C0MoERR<(02RE
CMRRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRbDV0C$bRR:=O#DN#RVb5RD,VNDF0E_OC_O	CFsss
2;RRRRRVRsbb0$C=R:RNOD#b#VR,5sRFVDNO0_E	CO_sCsF;s2
RRRR8CMR;HV
RRRRRHV5bDV0C$bRM=RCxo_CRsFFDsRV$b0b=CRR#bF_sxCFN2RMR8
RRRRRV5sbb0$CRR=M_CoxFCsRRFss0Vb$RbC=FRb#C_xsRF20MEC
RRRRHRR#J_CkRND:'=R4
';RRRRCCD#
RRRRDRRsHC#x:CR=CRs#CHxRs5NoRRRRRRRRRRRRR=>DR,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>VNDF0C_8MlFsNxDHCR,
RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>DRVF_N08FCMsDlNH2xC;R
RRRRRs#sCHRxC:s=RCx#HCNR5sRoRRRRRRRRRR>R=R
s,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RFVDN80_CsMFlHNDx
C,RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=V>RD0FN_M8CFNslDCHx2R;
RRRRR_H#CNJkD=R:R_0F#PkD5CDs#CHx2=R?R_0F#PkD5Css#CHx2R;
RCRRMH8RVR;
RHRRVVR5D0FN_COEOC	_sssF2ER0CRM
RRRRRRHV5bDV0C$bRM=RNFMRsVRDbb0$CRR=JCkH0N_MMsRF
RRRRRRRRsRRV$b0b=CRRMMNRRFss0Vb$RbC=kRJH_C0M2NMRC0EMR
RRRRRR#RH_FkMss8CC:8R=4R''R;
RRRRR#CDCR
RRRRRR#RH_FkMss8CC:8R=jR''R;
RRRRR8CMR;HV
RRRR#CDCR
RRRRRHk#_M8FsC8sCRR:=';j'
RRRR8CMR;HV
RRRR0sCkRsMMRF05_H#CNJkDMRN8FRM0#RH_FkMss8CC;82
CRRMV8Rk0MOHRFM"=?/"
;
RkRVMHO0F"MR?R>"5Rp,)RR:z h)1emp V7_D0FN2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=-MlHC'5DD,FIRDs'F;I2
RRRRsPNHDNLCFRVk8M8NR#ERRRRRA:Rm mpq:hR=NRVD;#C
LRRCMoH
RRRRRHV5NVsOF0HMH_I8R0E=RRjFDsR'MDCoR0E<RR(FssR'MDCoR0E<2R(RC0EMR
RRRRRskC0s'MRX
';RRRRCCD#
RRRRVRRFHsRRRHMpN'sMRoCDbFF
RRRRRRRRRHVp25HR'=R-0'RE
CMRRRRRRRRRFRVk8M8NR#E:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRVRRFHsRRRHM)N'sMRoCDbFF
RRRRRRRRRHV)25HR'=R-0'RE
CMRRRRRRRRRFRVk8M8NR#E:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRHRRVFRVk8M8NR#E0MEC
RRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRRRRR&""R"?">":-R''FRVkRM8HOMRFNlbs#CR0MsHoR"
RRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRR0sCkRsM';X'
RRRRCRRDV#HR_H#G25DRRFsHG#_5Rs20MEC
RRRRRRRR0sCkRsM';X'
RRRRCRRDV#HR>DRR0sRE
CMRRRRRRRRskC0s'MR4
';RRRRRDRC#RC
RRRRRsRRCs0kMjR''R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMV8Rk0MOHRFM""?>;R

RMVkOF0HM?R">R="5Rp,)RR:z h)1emp V7_D0FN2CRs0MksR71a_mzptRQBHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=-MlHC'5DD,FIRDs'F;I2
RRRRsPNHDNLCFRVk8M8NR#ERRRRRA:Rm mpq:hR=NRVD;#C
LRRCMoH
RRRRRHV5NVsOF0HMH_I8R0E=RRjFDsR'MDCoR0E<RR(FssR'MDCoR0E<2R(RC0EMR
RRRRRskC0s'MRX
';RRRRCCD#
RRRRVRRFHsRRRHMpN'sMRoCDbFF
RRRRRRRRRHVp25HR'=R-0'RE
CMRRRRRRRRRFRVk8M8NR#E:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRVRRFHsRRRHM)N'sMRoCDbFF
RRRRRRRRRHV)25HR'=R-0'RE
CMRRRRRRRRRFRVk8M8NR#E:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRHRRVFRVk8M8NR#E0MEC
RRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRRRRR&""R"?">="':R-V'RF8kMRRHMObFlNRsC#H0sM
o"RRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRCRs0MksR''X;R
RRRRRCHD#V#RH_DG52sRFR_H#G25sRC0EMR
RRRRRRCRs0MksR''X;R
RRRRRCHD#VRRD>s=RRC0EMR
RRRRRRCRs0MksR''4;R
RRRRRCCD#
RRRRRRRR0sCkRsM';j'
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R">;="
R
RVOkM0MHFR<"?"pR5,RR):hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;
RPRRNNsHLRDCVMFk8#8NERRRR:RRRmAmph qRR:=V#NDCR;
RoLCHRM
RHRRVVR5s0NOH_FMI0H8ERR=jsRFRDD'C0MoERR<(sRFRDs'C0MoERR<(02RE
CMRRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRsVFRHHRM'RpsoNMCFRDFRb
RRRRRHRRV5RpH=2RR''-RC0EMR
RRRRRRRRRVMFk8#8NE=R:Rk0sCR;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRVMFk8#8NE=R:Rk0sCR;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRRHVVMFk8#8NEER0CRM
RRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCR
RRRRRRRRR&RR""<"?"R":'R-'VMFk8MRHRlOFbCNsRs#0H"Mo
RRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRsRRCs0kMXR''R;
RRRRR#CDHHVR#5_GDF2Rs#RH_sG52ER0CRM
RRRRRsRRCs0kMXR''R;
RRRRR#CDHDVRRs<RRC0EMR
RRRRRRCRs0MksR''4;R
RRRRRCCD#
RRRRRRRR0sCkRsM';j'
RRRRCRRMH8RVR;
RCRRMH8RVR;
R8CMRMVkOF0HM?R"<
";
VRRk0MOHRFM"=?<"pR5,RR):hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=lR-H5MCDF'DIs,R'IDF2R;
RPRRNNsHLRDCVMFk8#8NERRRR:RRRmAmph qRR:=V#NDCR;
RoLCHRM
RHRRVVR5s0NOH_FMI0H8ERR=jsRFRDD'C0MoERR<(sRFRDs'C0MoERR<(02RE
CMRRRRRCRs0MksR''X;R
RRDRC#RC
RRRRRsVFRHHRM'RpsoNMCFRDFRb
RRRRRHRRV5RpH=2RR''-RC0EMR
RRRRRRRRRVMFk8#8NE=R:Rk0sCR;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRsVFRHHRM'R)soNMCFRDFRb
RRRRRHRRV5R)H=2RR''-RC0EMR
RRRRRRRRRVMFk8#8NE=R:Rk0sCR;
RRRRRCRRMH8RVR;
RRRRR8CMRFDFbR;
RRRRRRHVVMFk8#8NEER0CRM
RRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCR
RRRRRRRRR&RR""<"?=:""R''-RkVFMH8RMFROlsbNC0R#soHM"R
RRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRskC0s'MRX
';RRRRRDRC#RHVHG#_5RD2FHsR#5_Gs02RE
CMRRRRRRRRskC0s'MRX
';RRRRRDRC#RHVD=R<R0sRE
CMRRRRRRRRskC0s'MR4
';RRRRRDRC#RC
RRRRRsRRCs0kMjR''R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMV8Rk0MOHRFM"=?<"
;
RkRVMHO0F#MR0l8_NE0OR,5pR:)RR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRRRHV5Ep'HRoE='R)EEHoR8NMRDp'F=IRRD)'FRI20MEC
RRRRsRRCs0kM0R#8N_l05OE0#F_k5DPpR2,0#F_k5DP);22
RRRR#CDCR
RRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_MlRC
RRRRR&RRRa"17q_va:B]R)p'q htRR/=)q')h,t R0sCkHsMMwoRq p1"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRDVN#
C;RRRRCRM8H
V;RMRC8kRVMHO0F#MR0l8_NE0O;R

RMVkOF0HMHRVMs8_H0oEl0F#Rs5NoRR:z h)1emp V7_D0FN;RR$:aR17p_zmBtQ2CRs0MksRaQh )t R
H#RCRLo
HMRRRRV_FsDbFFRV:RFHsRRRHMN'sosCCPs_#CsoNMCFRDFRb
RRRRRRHVN5soH?2R=RR$0MEC
RRRRRRRR0sCkRsMHR;
RRRRR8CMR;HV
RRRR8CMRFDFbR;
RsRRCs0kMsRNoH'Eo4E+;RRRRRRRRRRRRRRRR-RR-CRs0MksR0FkRRFVLMFk8'#REEHo
CRRMV8Rk0MOHRFMV8HM_osHEF0l#
0;
VRRk0MOHRFMV8HM_VDC0#lF0NR5s:oRR)zh p1me_ 7VNDF0$;RR1:Raz7_pQmtBs2RCs0kMhRQa  t)#RH
LRRCMoH
RRRRsVF_FDFbRR:VRFsHMRHRoNs'MsNoDCRF
FbRRRRRVRHRoNs5RH2?$=RRC0EMR
RRRRRRCRs0MksR
H;RRRRRMRC8VRH;R
RRMRC8FRDF
b;RRRRskC0sNMRsDo'F4I-;RRRRRRRRRRRRRRRRRRR-s-RCs0kMkRF0VRFRkLFMR8#'IDF
CRRMV8Rk0MOHRFMV8HM_VDC0#lF0
;
R-R-RCaE#FCRPsCsHR8C0REC8NCVk#D0RsVFRC0ERlOFbCNsRCFbsFN0s
#3RkRVMHO0F"MR=5"RDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMJRC5RD,s
2;RMRC8kRVMHO0F"MR=
";
VRRk0MOHRFM""/=R,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMMDC5,2Rs;R
RCRM8VOkM0MHFR="/"
;
RkRVMHO0F"MR>R="5RD,sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0soMRC,5DR;s2
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"RDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm RqhHR#
RoLCHRM
RsRRCs0kMCRD5RD,s
2;RMRC8kRVMHO0F"MR<;="
R
RVOkM0MHFR"">R,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
LRRCMoH
RRRR0sCkRsMoD05,2Rs;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""DR5,RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpqHhR#R
RLHCoMR
RRCRs0MksR5D0Ds,R2R;
R8CMRMVkOF0HM<R""
;
R-R-RsbkbCF#:NRlGkHllVRFRF0IRlMkL#CsRP5FCHss8RC#8NCVk2D0
VRRk0MOHRFMlHNGlRkl5R
RR,RpR:)RR)zh p1me_ 7VNDF0R2
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0ERRR:hzqa)Rqp:-=RlCHM5DD'FRI,sF'DIR2;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0GRCbCFMMI0_HE80R:RRRahqzp)qRR:=lHNGl5klDH'EoRE,sH'Eo;E2R-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHNDDCRsHC#xRC,s#sCHRxC:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RCRLo
HMRRRRH5VR5Dp'C0MoERR<4F2Rs)R5'MDCoR0E<2R42ER0CsMRCs0kMqRhw
u;RRRRCRM8H
V;RRRRD#sCHRxC:s=RCx#HCDR5,GRCbCFMMI0_HE80,sRVNHO0FIM_HE802R;
RsRRsHC#x:CR=CRs#CHxR,5sRbCGFMMC0H_I8,0ERNVsOF0HMH_I820E;R
RRVRHRCDs#CHxRs>RsHC#x0CRERCMskC0sDMRsHC#x
C;RRRRCCD#R0sCkRsMs#sCH;xC
RRRR8CMR;HV
CRRMV8Rk0MOHRFMlHNGl;kl
R
RVOkM0MHFRMlHHllkRR5
RpRR,RR):hRz)m 1p7e _FVDN
02RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0sRVNHO0FIM_HE80R:RRRahqzp)qRR:=-MlHC'5DD,FIRDs'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERRR:qRhaqz)p=R:RGlNHllk5ED'H,oEREs'H2oE;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RPRRNNsHLRDCD#sCH,xCRCss#CHxRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
LRRCMoH
RRRRRHV5'5pDoCM0<ERRR42F5sR)C'DMEo0R4<R202RERCMskC0shMRq;wu
RRRR8CMR;HV
RRRRCDs#CHxRR:=sHC#x5CRDC,RGMbFC_M0I0H8EV,Rs0NOH_FMI0H8E
2;RRRRs#sCHRxC:s=RCx#HCsR5,GRCbCFMMI0_HE80,sRVNHO0FIM_HE802R;
RHRRVsRDCx#HCRR>s#sCHRxC0MECR0sCkRsMs#sCH;xC
RRRR#CDCCRs0MksRCDs#CHx;R
RRMRC8VRH;R
RCRM8VOkM0MHFRMlHHllk;R

R----------------------------------------------------------------------------R-
RR--OPFMCHs#FVMRk0MOH#FM
-RR----------------------------------------------------------------------------
R
R-B-RFCMPsR0#NDRVFHN0MboRF0HMRlMkLRCsFFVRMVCRFNsl0MRH0NFRMEF0CVsRFNsl0R
RVOkM0MHFR#sCHRxC5R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRRRRRRRR--wNDF0oHMRHbFMH0RM0bk
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azqRpRR=R:RFVDNC0_GMbFC_M0I0H8ER;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)pRRRRR:=VNDF0s_VNHO0FIM_HE80;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0sMFk80_#$RDCR:RRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsFRsRRRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;Fs
RRRRMOF#M0N0CR8MlFsNxDHCM_HRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC;RR--zR#CQ   R0CGCCM88uRw
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRFROMN#0MH0RMs_VNHO0FIM_HE80Rh:Rq)azq:pR=NR-sDo'FRI;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0MRH_bCGFMMC0H_I8R0E:qRhaqz)p=R:RoNs'oEHER;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRPHNsNCLDR#sCkRD0RRRRRRRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-CRs#0kDRDPNkRC
RPRRNNsHLRDCV$b0bRCRRRRRRRRRRRR:PHND8b_V#00NCR;
RPRRNNsHLRDCCFGbMM_HRRRRRRRRRRR:1hQt 57RHCM_GMbFC_M0I0H8ER-48MFI0jFR2R;
RPRRNNsHLRDCVOsN0M_HRRRRRRRRRRR:zQh1t7h RM5H_NVsOF0HMH_I8R0E8MFI0jFR2R;
RPRRNNsHLRDCsMFk8RRRRRRRRRRRRRR:Apmm ;qh
RRRRsPNHDNLCGRCb_FMFRk0RRRRRRRR:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2Rj;-RR-kRF00bkRNVsOR0
RPRRNNsHLRDCVOsN0k_F0RRRRRRRRRR:zQh1t7h Rs5VNHO0FIM_HE80RI8FMR0FjR2;RR--Fbk0kV0Rs0NO
RRRRsPNHDNLCNRb#k#oNRs8RRRRRRRR:qRhaqz)pR;
RoLCHRM
RVRRbb0$C=R:RNOD#b#V5oNs,EROC_O	CFsss
2;RRRRH5VR50Vb$RbC=FRb#C_8MlFsNFDRsbRV0C$bRM=RC8o_CsMFl2NDR8NMRM8CFNslDCHx_
HMRRRRRRRRNRM85_HMCFGbM0CM_8IH0<ERRbCGFMMC0H_I8
0ERRRRRRRRRRRRRRFsHVM_s0NOH_FMI0H8ERR<VOsN0MHF_8IH02E2
RRRRFRRsMRH_bCGFMMC0H_I8R0E>GRCbCFMMI0_HE80
RRRRFRRsMRH_NVsOF0HMH_I8R0E>sRVNHO0FIM_HE80RC0EMR
RRRRR-#-RHRxCskC8OF0HMR
RRRRRO#DN##ONCRR:OCN#R0Vb$RbCHR#
RRRRRIRRERCMHR#G=R>
RRRRRRRRR#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRRRRRIMECRMMNRJ|Rk0HC_MMNR
=>RRRRRRRRRCRs#0kDRR:=JMMNV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRCIEMFRb#M_HV>R=
RRRRRRRRsRRCD#k0=R:R#bF_VHMV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRIMECRoMC_VHMR
=>RRRRRRRRRCRs#0kDRR:=M_CoHVMVbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRIRRERCMb_F#xFCsRM|RCxo_CRsF=R>
RRRRRRRRR#sCkRD0:x=RCVsFbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0ER-RR-NRE0-CRjR
RRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRCIEM0RFE#CsR
=>RRRRRRRRRsRLC_N	MLklC5sR
RRRRRRRRRRRRoNsRRRRRRRRRR=>N,so
RRRRRRRRRRRR0Vb$RbRRRRRRR=>V$b0b
C,RRRRRRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDxHC_MR,
RRRRRRRRRVRRs0NORRRRR=RR>sRVN_O0H
M,RRRRRRRRRRRRCFGbMRRRRRRR=C>RGMbF_2HM;R
RRRRRRRRRHVVRs0NOH_FMI0H8ERR>HVM_s0NOH_FMI0H8EMRN8CR8MlFsNxDHCM_HRC0EMR
RRRRRRRRRR-R-RkYFRDFM$CRo0CREsHCRVFR$kNREPNCRRM8CFNslDMRHb
k0RRRRRRRRRRRRVOsN0k_F0=R:R05FE#CsRR=>'2j';RRRRRRRRRRRR-RR-NRb8HRI0xERC#sF
RRRRRRRRRRRRNVsOF0_k50RVOsN0MHF_8IH08ERF0IMFR
RRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E-MRH_NVsOF0HMH_I820ERR:=VOsN0M_H;R
RRRRRRRRRRCRs#0kDRR:=MlFsNxDHC
R5RRRRRRRRRRRRRsRVNRO0RRRRRRRRRR=>VOsN0k_F0R,
RRRRRRRRRRRRRbCGFRMRRRRRRRRR=C>RGMbF_,HM
RRRRRRRRRRRR#RRHRoMRRRRRRRRR>R=RoNs5oNs'oEHE
2,RRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRMNoksR8RRRRRR=RR>2Rj;R
RRRRRRRRRCCD#
RRRRRRRRRRRR#sCkRD0:M=RFNslDCHxRR5
RRRRRRRRRRRRRNVsOR0RRRRRRRRR=V>Rs0NO_,HM
RRRRRRRRRRRRCRRGMbFRRRRRRRRR>R=RbCGFHM_MR,
RRRRRRRRRRRRRo#HMRRRRRRRRRRR=N>RsNo5sEo'H2oE,R
RRRRRRRRRRRRRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx
C,RRRRRRRRRRRRRoRMk8NsRRRRRRRRRR=>HVM_s0NOH_FMI0H8ERR-VOsN0MHF_8IH0;E2
RRRRRRRRCRRMH8RVR;
RRRRR8CMR#ONCDRONO##N;#C
RRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--#CHxROHMs#CNCsRFRC0ERl#NCHR#xRC
RRRRRRHVCFGbM0CM_8IH0>ERR_HMCFGbM0CM_8IH00ERE
CMRRRRRRRRCFGbMM_HRR:=1hQt N75s5oRHCM_GMbFC_M0I0H8ER-48MFI0jFR2
2;RRRRRRRRHVVRbb0$CRR=b_F#xFCsRRFsV$b0b=CRRoMC_sxCFER0CRM
RRRRRRRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>jR''
2;RRRRRRRRCHD#VGRCb_FMH=MRRR-40MECRRRRRRRR-H-RMFVRsNRMM#R5E0Fs#kRF0EROC_O	CFsssR2
RRRRRRRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>4R''
2;RRRRRRRRCCD#
RRRRRRRR-RR-MRHP0CsRb0FRaAQ
RRRRRRRRCRRGMbF_5HMCFGbMM_H'oEHER2RRR:=MRF0CFGbMM_H5bCGFHM_MH'Eo;E2
RRRRRRRRCRRGMbF_0FkRR:=sHC#x5CRCFGbMM_H,GRCb_FMF'k0DoCM0;E2R-R-Ro#HMRC8CNGbMR8
RRRRRRRRRR--wbDHRRH0L	NO3R
RRRRRRRRRCFGbMk_F0G5Cb_FMF'k0EEHo2=R:R0MFRbCGFFM_kC05GMbF_0Fk'oEHE
2;RRRRRRRRRCRs#0kDRG5CbCFMMI0_HE80-84RF0IMF2RjRR:=z h)1emp V7_D0FN5bCGFFM_k;02
RRRRRRRR8CMR;HV
RRRRRRRR#sCkRD05bCGFMMC0H_I820ERR:=NRso5_HMCFGbM0CM_8IH0;E2RRRRRR--#MHo
RRRRCRRDR#CRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--CFGbM0CM_8IH0=ERR_HMCFGbM0CM_8IH0RE
RRRRRsRRCD#k0CR5GMbFC_M0I0H8EFR8IFM0RRj2:N=Rs5oRHCM_GMbFC_M0I0H8EFR8IFM0R;j2
RRRRCRRMH8RVR;
RRRRRRHVVOsN0MHF_8IH0>ERR_HMVOsN0MHF_8IH00ERE
CMRRRRRRRRskC#D50R-84RF0IMFVR-s0NOH_FMI0H8E:2R=FR50sEC#>R=R''j2R;R-x-RC#sF
RRRRRRRR#sCkRD05R-48MFI0-FRHVM_s0NOH_FMI0H8E:2R=R
RRRRRRRRRNRso5R-48MFI0-FRHVM_s0NOH_FMI0H8E
2;RRRRRDRC#RCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-V-Rs0NOH_FMI0H8ERR=HVM_sHNO0_FMI0H8ER
RRRRRRCRs#0kDR45-RI8FMR0F-NVsOF0HMH_I820ER
:=RRRRRRRRRsRNo-R54FR8IFM0RM-H_NVsOF0HMH_I820E;R
RRRRRCRM8H
V;RRRRCRM8H
V;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMCRs#CHx;R

RMVkOF0HMCRs#CHxRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRRRR:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFsR:RRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDxHC_MRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0#R5H_xCs'C#D0CVRI8FMR0F#CHx_#sC'osHE;02
LRRCMoH
RRRRRHV5#sCk'D0DoCM0<ERRR420MEC
RRRRsRRCs0kMCRs#0kD;R
RRDRC#RC
RRRRR#sCkRD0:s=RCx#HCNR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRORRE	CO_sCsFRsRR>R=RCOEOC	_sssF,R
RRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH_xCH
M,RRRRRRRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHC
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFMsHC#x
C;
VRRk0MOHRFM0VF_D0FNd5.R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRCOEOC	_sssFRRRR:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;
RORRF0M#NRM08FCMsDlNH_xCH:MRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx;-RR-#RzC RQ C RGM0C8RC8wRu
RORRF0M#NRM08FCMsDlNHRxCR:RRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDN.0dR
H#RCRLo
HMRRRRskC0ssMRCx#HCNR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=V>RD0FNdE.'H,oE
RRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>VR-D0FNdD.'F
I,RRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRCOEOC	_sssFRRRR=O>RE	CO_sCsF
s,RRRRRRRRRRRRRRRRR8RRCsMFlHNDxHC_M>R=RM8CFNslDCHx_,HM
RRRRRRRRRRRRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHC
2;RMRC8kRVMHO0F0MRFD_VFdN0.
;
RkRVMHO0F0MRFD_VFnN0c
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRRRR:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFsR:RRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDxHC_MRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0RncHR#
RoLCHRM
RsRRCs0kMCRs#CHxRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>DRVFnN0cH'Eo
E,RRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RD-VFnN0cF'DIR,
RRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRROOEC	s_CsRFsR=RR>EROC_O	CFsssR,
RRRRRRRRRRRRRRRRRCR8MlFsNxDHCM_HRR=>8FCMsDlNH_xCH
M,RRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
R8CMRMVkOF0HMFR0_FVDNc0n;R

RMVkOF0HMFR0_FVDN.04U
R5RRRRNRsoRRRRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRRRR:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFsR:RRRmAmph qRRRR:V=RD0FN_COEOC	_sssF;R
RRFROMN#0M80RCsMFlHNDxHC_MRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH;xCR-R-RCz#R Q  GRC08CMCw8RuR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCz#R Q  GRC08CMCw8RuR
RRCRs0MksR)zh p1me_ 7VNDF0U4.R
H#RCRLo
HMRRRRskC0ssMRCx#HCNR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=V>RD0FN4'.UEEHo,R
RRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=->RVNDF0U4.'IDF,R
RRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRORRE	CO_sCsFRsRR>R=RCOEOC	_sssF,R
RRRRRRRRRRRRRRRRRRM8CFNslDCHx_RHM=8>RCsMFlHNDxHC_MR,
RRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RCRM8VOkM0MHFR_0FVNDF0U4.;R

RR--0VF_D0FNRC5)N
D2R-R-Rb0$HDONDM$RF10R$EM0Cx#HNCLDRDkMCR##0RECHkMb0#RHRONRF0M#N3M0
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRRq) pR;
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLCsRNoC_sNRDRR):R ;qpRRRRRRRRRR--)DCNRsPC#MHFRRFVNksol0CM
RRRRsPNHDNLCNRPDVH8bRRRRL:RF8kMN_s$0C$b;RRRR-RR-ERBCRO	VRFsPHND8CRs#0kD#R
RRNRPsLHNDCCRGRbRRRRRRRR:Q hat; )RRRRR-R-R0QMCsoCRsPC#MHFRRFVCFGbM0CM
RRRRsPNHDNLCGRCbRFMRRRRRz:Rht1QhR 75bCGFMMC0H_I8R0E-RR48MFI0jFR2R;
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-MRz#MHoCP8RCHs#FFMRVGRCbR3
RORRF0M#NRM0CFGbMN_L#:CRRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0RRj2:R=
RRRRRMoC_bCGFLM_N5#CCFGbM0CM_8IH0;E2R-RR-GRCbCFMMF0RVCV#0R
RRNRPsLHNDVCRs0NORRRRRz:Rht1QhR 75NVsOF0HMH_I8-0E4FR8IFM0R;j2
RRRRsPNHDNLCsRVNRORRRRR: R)qRp;RRRRRRRRRR--)DCNRsPC#MHFRRFVVOsN0MHF
RRRRMOF#M0N0FRskVM8sRNO: R)q:pR=3R.j*R*R.5-RV-Rs0NO'oEHER2;RR--k8#CRsVFRksFMM8HoR
RRNRPsLHNDsCRF8kMRRRRRA:Rm mpqRh;RRRRR-R-RR0FsMFk8sRFR0MFRR0FsMFk8R
RLHCoMR
RRCRs#0kDR:RR=FR50sEC#>R=R''j2R;
RNRRsso_CRND:N=Rs
o;RRRRHNVRsso_CRND<3RjjER0CRM
RRRRR#sCkRD05bCGFMMC0H_I820ERR:=';4'
RRRRNRRsso_CRNDRRRRRRRRRRRRR:RR=RR-N_sosDCN;-RR-NRv	HCR0FRb#HH0P
C3RRRRCCD#
RRRRsRRCD#k0CR5GMbFC_M0I0H8E:2R=jR''R;
RCRRMH8RVR;
R0RRC_#0LMFk8$NsRs5NoRRRRRRRRRRRRR=>N_sosDCN,R
RRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0
E,RRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx,R
RRRRRRRRRRRRRRRRRR$L0bRCRRRRRRRRR=P>RN8DHV
b,RRRRRRRRRRRRRRRRRDRRFHo.RRRRRRRRR>R=RbCG2R;
RHRRVNRPDVH8bRR=xFCsRC0EMR
RRRRRskC0ssMRCD#k0R;RRRRRRRRRRRRRRRRRR-R-R#)CkRD0H0MHHHNDxRC80"FRj
"3RRRRCHD#VNRPDVH8bRR=HHMVM$H0RC0EMR
RRRRRskC#D50RCFGbM0CM_8IH0-ERR84RF0IMF2RjRR:=5EF0CRs#='>R4;'2R-R-Rb GFMMC0DRND4R""R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-R-R0sCkRsMHHMVM$H03R
RRRRRskC0ssMRCD#k0R;
RCRRD
#CRRRRRVRHRDPNHb8VR8=RCsMFlRND0MECRRRRRRRR- -RGMbFCRM0IDHDRV8CN0kDRR0F"3j"
RRRRRRRRbCGF:MR=FR50sEC#>R=R''j2R;
RRRRRVRRsRNORR:=N_sosDCNR5*R.R3j*5*R0HF_Mo0CCCs5GMbF_#LNC42-2
2;RRRRRDRC#RCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-h-RkClLsCRD#0#RERNM4"3RMlFsNRD"MLklCRs
RRRRRCRRGMbFRRRR:z=Rht1QhR 75_0F#MHoC58RC-Gb4C,RGMbFC_M0I0H8E;22
RRRRRRRRbCGFCM5GMbFC_M0I0H8E2-4RR:=MRF0CFGbMG5CbCFMMI0_HE80-;42
RRRRRRRRNVsORRRR=R:Rs5NoC_sN/DRRj.3RR**C2GbR4-R3Rj;RR--hLklCDsRCR##0MENR
43RRRRRMRC8VRH;R
RRRRRVRFsHMRHR0jRFsRVN'O0EEHoRFDFbR
RRRRRRVRHRNVsO=R>Rj.3RR**5R-4-2RHRC0EMR
RRRRRRRRRVOsN0VR5s0NO'oEHERR-H:2R=4R''R;
RRRRRRRRRNVsORRRRRRRRRRRRRRRRRRR:V=RsRNO-3R.j*R*R45-RH-R2R;
RRRRRCRRD
#CRRRRRRRRRsRVNRO05NVsOE0'HRoE-2RHRR:=';j'
RRRRRRRR8CMR;HV
RRRRCRRMD8RF;Fb
RRRRsRRF8kMRR:=V#NDCR;
RRRRR#ONCFRsk_M8#D0$C#RH
RRRRRRRRCIEMFRsk_M8MsCNCR#0=R>
RRRRRRRRRRHVVOsNRs>RF8kMVOsNRRFs5s5VN=ORRksFMs8VNRO2NRM8VOsN025jR'=R4R'20MEC
RRRRRRRRRRRRksFM:8R=sR0k
C;RRRRRRRRRMRC8VRH;R
RRRRRRERICsMRF8kM_VHMR
=>RRRRRRRRRVRHRNVsO=R/Rjj3R8NMR#sCk5D0CFGbM0CM_8IH0RE2=jR''ER0CRM
RRRRRRRRRsRRF8kMRR:=0Csk;R
RRRRRRRRRCRM8H
V;RRRRRRRRIMECRksFMM8_CMoHV>R=
RRRRRRRRHRRVsRVN/OR=3RjjMRN8CRs#0kD5bCGFMMC0H_I820ER'=R40'RE
CMRRRRRRRRRRRRsMFk8=R:Rk0sCR;
RRRRRRRRR8CMR;HV
RRRRRRRRCIEM0RFE#CsR
=>RRRRRRRRRkRMDRD;RRRRRRRRRRRRRRRRRRRRRRRR-8-RF0M'RksFMR8
RRRRR8CMR#ONCR;
RRRRRRHV5ksFMR820MEC
RRRRRRRRRHVN5M8VOsN0=2RR''4RC0EMRRRRRRRRR--VOsN0MHFRRH#NRDD"
4"RRRRRRRRRGRCbRFM:C=RGMbFR4+R;R
RRRRRRRRRVOsN0=R:R05FE#CsRR=>'2j';R
RRRRRRDRC#RC
RRRRRRRRRNVsO:0R=sRVNRO0+;R4
RRRRRRRR8CMR;HV
RRRRCRRMH8RVR;
RRRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:z=Rh1) m pe7D_VF5N0CFGbM
2;RRRRRCRs#0kDR45-RI8FMR0F-NVsOF0HMH_I820ERR:=z h)1emp V7_D0FN5NVsO;02
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-R_0FVNDF0QR5Mo0CC
s2RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:Q hat; )
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azqRpRR=R:RFVDNC0_GMbFC_M0I0H8ER;R-D-RC0MoEVRFRRwuFbk0kC0RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)pRRRRR:=VNDF0s_VNHO0FIM_HE80;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0sMFk80_#$RDCR:RRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D2-RR-FRskHM8MFoRbF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#DR0RR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RPRRNNsHLRDCN_soHRM0R:RRRahqzp)q;RRRR-RR-NRh0NksDCRPsF#HMVRFRoNskMlC0R
RRNRPsLHNDCCRGMbFRRRRRRR:1hQt 57RCFGbM0CM_8IH04E-RI8FMR0Fj
2;RRRRPHNsNCLDRbCG0RlbRRRR:QR1t7h RG5CbCFMMI0_HE80-84RF0IMF2Rj;R
RR-R-R#zMHCoM8CRPsF#HMVRFRbCG3R
RRFROMN#0MC0RGMbF_#LNCRR:1hQt 57RCFGbM0CM_8IH04E-RI8FMR0Fj:2R=R
RRRRRo_CMCFGbMN_L#CC5GMbFC_M0I0H8ER2;R-R-RbCGFMMC0VRFV0#C
RRRRsPNHDNLCsRVNRO0RRRR:hRz1hQt 57RVOsN0MHF_8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''j2R;
RPRRNNsHLRDCVOsN0b0lRRR:zQh1t7h Rs5VNHO0FIM_HE80-84RF0IMF2Rj;R
RRNRPsLHNDsCRF8kMRRRRRA:Rm mpq
h;RRRRPHNsNCLDRH#EVR0RR:RRRahqzp)q;R
RRNRPsLHND#CRE0HVsRRRRh:Rq)azq
p;RRRRPHNsNCLDRksFMs8VN:ORRahqzp)q;RRRRRRR-k-R#RC8HsMRF8kMH
MoRCRLo
HMRRRRHNVRs<oRR0jRE
CMRRRRRCRs#0kDRG5CbCFMMI0_HE802=R:R''4;R
RRRRRN_soHRM0RRRRRRRRRRRRRRRR:-=RN;soR-R-R	vNC0RHR#bFHP0HCR3
RCRRD
#CRRRRRCRs#0kDRG5CbCFMMI0_HE802=R:R''j;R
RRRRRN_soHRM0RRRRRRRRRRRRRRRR:N=Rs
o;RRRRCRM8H
V;RRRRHNVRsHo_M=0RR0jRE
CMRRRRRCRs#0kDRR:=xFCsV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRR#CDCR
RRRRR-Q-RVER0CkRMlsLCRRH#DoNsC0sRERNMIOCRNsMRCCbs#0CMRRHM0#EHRlMkLRCs#0$#CRl
RRRRRR--IMCRCRC80sFRCs0kMMRHVHHM0
$3RRRRRER#HRV0:D=RF5o.N_soH2M0;R
RRRRRH#VRE0HVR0>RFM_H0CCosG5Cb_FMLCN#2ER0CRM
RRRRR-RR-FRIsRs$NkLF0MRHVHHM0R$
RRRRRHRRVCRs#0kDRG5CbCFMMI0_HE802RR='Rj'0MEC
RRRRRRRRsRRCD#k0=R:R#bF_VHMV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRCCD#
RRRRRRRR-RR-CRs0MksRoMCNP0HCMRHVHHM0
$3RRRRRRRRRCRs#0kDRR:=M_CoHVMVbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRCRRMH8RVR;
RRRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-FRhsDlNRlMkLRCs5MON'L0RCCR8MlFsN
D2RRRRRRRR-B-RFklb0 CRGMbFC
M0RRRRRRRRCFGbMRRR:0=RFH_#o8MCRE5#H-V04C,RGMbF'MDCo20E;-RR-FRb#HH0PVCRs0NOH3FM
RRRRRRRRR--BbFlkR0CwOsN0MHF
RRRRRRRRoNs_0HMRR:=N_soHRM0-*R.*H#EVR0;RR--10kLs0NORVFVRC0ERj43
RRRRRRRRH#EVR0sRR:=#VEH0R;
RRRRRVRRFQsRRRHMVOsN0H'Eo8ERF0IMFNRlGkHllVR5s0NO'oEHERR-#VEH0RR+4j,R2FRDFRb
RRRRRRRRRH#EVR0s:#=RE0HVsRR-4R;
RRRRRRRRRRHV5oNs_0HMRR>=.#**E0HVs02RE
CMRRRRRRRRRRRRN_soHRM0RR:=N_soHRM0-*R.*H#EV;0s
RRRRRRRRRRRRNVsOQ052=R:R''4;R
RRRRRRRRRCCD#
RRRRRRRRRRRRNVsOQ052=R:R''j;R
RRRRRRRRRCRM8H
V;RRRRRRRRCRM8DbFF;R
RRRRRR-R-Rk)FMM8HoFRskM0HCR
RRRRRRFRskRM8:V=RNCD#;R
RRRRRRVRHRoNs_0HMRj>RRC0EMR
RRRRRRRRRsMFk8NVsO=R:R*.*5H#EV-0s4
2;RRRRRRRRRNRO#sCRF8kM_$#0DHCR#R
RRRRRRRRRRERICsMRF8kM_NMCs0C#R
=>RRRRRRRRRRRRRVRHRoNs_0HMRs>RF8kMVOsNR
FsRRRRRRRRRRRRRRRR5s5NoM_H0RR=sMFk8NVsON2RMV8Rs0NO5Rj2=4R''02RE
CMRRRRRRRRRRRRRRRRsMFk8=R:Rk0sCR;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRCIEMFRsk_M8HRMV=R>
RRRRRRRRRRRRRRHVN_soHRM0/j=RR8NMR#sCkRD05bCGFMMC0H_I820ER'=Rj0'RE
CMRRRRRRRRRRRRRRRRsMFk8=R:Rk0sCR;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRCIEMFRsk_M8MHCoM=VR>R
RRRRRRRRRRRRRHNVRsHo_M/0R=RRjNRM8skC#D50RCFGbM0CM_8IH0RE2=4R''ER0CRM
RRRRRRRRRRRRRsRRF8kMRR:=0Csk;R
RRRRRRRRRRRRRCRM8H
V;RRRRRRRRRRRRIMECREF0CRs#=R>
RRRRRRRRRRRRRDMkDR;
RRRRRRRRR8CMR#ONCR;
RRRRRCRRMH8RVR;
RRRRRHRRVFRskRM80MEC
RRRRRRRRVRRbF_sk5M8VOsN0M_HR>R=RNVsO
0,RRRRRRRRRRRRRRRRRCRRGMbF_RHMRR=>CFGbMR,
RRRRRRRRRRRRRRRRRsRVN_O0FRk0=V>Rs0NO0,lb
RRRRRRRRRRRRRRRRRRRCFGbMk_F0>R=RbCG02lb;R
RRRRRRRRRVOsN0=R:RNVsOl00bR;
RRRRRRRRRbCGF:MR=GRCbb0l;R
RRRRRRMRC8VRH;R
RRRRRR-R-R0ukRC0ERlMkLRCs0CFo0sECR8NMR0sCk
sMRRRRRRRRCFGbMG5CbCFMMI0_HE80-R42RRRRRRRRR:RR=FRM0GRCb5FMCFGbM0CM_8IH04E-2R;
RRRRRsRRCD#k0CR5GMbFC_M0I0H8ER-48MFI0jFR2=R:R)zh p1me_ 7VNDF0G5Cb2FM;R
RRRRRRCRs#0kDR45-RI8FMR0F-NVsOF0HMH_I820ERR:=z h)1emp V7_D0FN5NVsO;02
RRRRCRRMH8RVR;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-R_0FVNDF0kR5Mo#HM2C8
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR1zhQ th7R;
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC2RR--sMFk8oHMR0FbH
FMRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RORRF0M#NRM0q_)tpa wRQ:Rhta  :)R=)RqtC'DMEo0-
4;RRRRNNDH#qRX)RtRRRRRRRR:zQh1t7h 5tq)_wp aFR8IFM0RRj2Hq#R)
t;RRRRPHNsNCLDRs#NoRRRRRR:1hQt 57Rq_)tpa w+84RF0IMF2Rj;-RR-HR#o8MCRsPC#MHFRRFVN
soRCRLo
HMRRRRHNVRsDo'C0MoERR<4ER0CRM
RRRRR0sCkRsMhuqw;R
RRMRC8VRH;R
RRNR#s5oRXtq)'MsNoRC2:1=RQ th7XR5q2)t;R
RRNR#s5oR#oNs'oEHER2R:'=Rj
';RRRRskC#D:0R=FR0_FVDN50RNRsoRRRRRRRRR=RR>NR#s
o,RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE80,R
RRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$C
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMFR0_FVDN
0;
-RR-FR0_FVDN50R#MHoC
82RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:1hQt 
7;RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)pRRRRR:=VNDF0G_CbCFMMI0_HE80;-RR-CRDMEo0RRFVwFuRkk0b0GRCbCFMMR0
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRRRR:V=RD0FN_NVsOF0HMH_I8;0ER-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$2DCR-R-RksFMM8HobRF0MHF
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RRRRRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RRFROMN#0Mq0R)pt_ RwaRRR:Q hatR ):q=R)Dt'C0MoE;-4
RRRRHNDNX#RqR)tRRRRRRRRR1:RQ th7)5qt _pw8aRF0IMF2RjRRH#q;)t
RRRRsPNHDNLCsRNoM_H0RRRRz:Rht1Qh5 7GoNs'MsNo;C2R-R-RN)CDCRPsF#HMVRFRoNskMlC0R
RRNRPsLHNDNCRs.oLRRRRRRR:zQh1t7h 5sGNoH'Eo.E/RI8FMR0FjR2;RR--D.FoRRFVHkMb0R
RRNRPsLHNDsCRCRGbRRRRRRR:1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj;R
RRNRPsLHNDCCRGRbRRRRRRRR:1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj;R
RR-R-Ro#HMRC8P#CsHRFMFCVRG
b3RRRRPHNsNCLDRbCGFRMRRRRR:hRz1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj;R
RR-R-R#zMHCoM8CRPsF#HMVRFRbCG3R
RRFROMN#0MC0RGMbF_#LNCRR:1hQt 57RCFGbM0CM_8IH04E-RI8FMR0Fj:2R=R
RRRRRo_CMCFGbMN_L#CC5GMbFC_M0I0H8ER2;R-R-RbCGFMMC0VRFV0#C
RRRRsPNHDNLCFRskRM8RA:Rm mpq
h;RRRRPHNsNCLDRNVsOR0R:hRz1hQt 57RVOsN0MHF_8IH04E-RI8FMR0Fj
2;RRRRPHNsNCLDRssVNRO0:hRz1hQt 57RVOsN0MHF_8IH04E-RI8FMR0Fj
2;RRRRPHNsNCLDRo#HMRRR:aR17p_zmBtQ;RRRRRRRR-R-Ro#HMHRL0R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR40MEC
RRRRsRRCs0kMqRhw
u;RRRRCRM8H
V;RRRRHQVR#R_X5sGNo02RE
CMRRRRRCRs#0kDRR:=5EF0CRs#='>RX;'2
RRRR#CDH5VRGoNsRj=R2ER0CRM
RRRRR#sCkRD0:x=RCVsFbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-h-RFNslDkRMlsLCRN5OMR'0L8CRCsMFl2ND
RRRR#RRHRoM:0=RFj_X4N5Gs5oRGoNs'oEHE;22
RRRRNRRsHo_M:0R=hRz1hQt N75L5#R0jF_4N5Gs2o22R;
RRRRRR--BbFlkR0C FGbM0CM
RRRRNRRs.oLRR:=0kF_Mo#HM5C8V8HM_VDC0#lF0s5NoM_H0',R4,'2RoNsLD.'C0MoER2;RR--p.Fo
RRRRHRRVsRNoRL.>hRz1hQt C75GMbF_#LNC02RE
CMRRRRRRRRskC#D:0R=FRb#M_HVRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRsRRCD#k0CR5GMbFC_M0I0H8E:2R=HR#o
M;RRRRRDRC#RC
RRRRRCRRGRbRR:RR=QR1t7h 5#sCH5xCNLso.C,RGDb'C0MoE;22
RRRRRRRRoNs_0HMRR:=#VEH0C_DV50RN_soH,M0RoNs_0HM'oEHEF-0_0HMCsoC5bCG2
2;RRRRRRRRH5VRN_soH'M0EEHoRV>Rs0NOH_FMI0H8E02RE
CMRRRRRRRRRsRVNRO0:N=RsHo_M50RN_soH'M0EEHo-84RF0IMFNR5sHo_ME0'H-oEVOsN0MHF_8IH02E2;R
RRRRRRRRRsMFk8=R:RCOEOs	_F8kMRR5
RRRRRRRRRVRRs0NO_RHMR=RR>sRVNRO05,j2
RRRRRRRRRRRRo#HMRRRRRRRRR=>#MHo,R
RRRRRRRRRRCRslMNH8RCsR>R=RoNs_0HM5s5NoM_H0H'EoVE-s0NOH_FMI0H8E2-4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8MFI0jFR2R,
RRRRRRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$C
2;RRRRRRRRRVRHRksFM08RE
CMRRRRRRRRRRRRVsb_F8kM5NVsOH0_M=RR>sRVN,O0
RRRRRRRRRRRRRRRRRRRRGRCb_FMHRMR=C>RG
b,RRRRRRRRRRRRRRRRRRRRRNVsOF0_k=0R>VRss0NO,R
RRRRRRRRRRRRRRRRRRCRRGMbF_0FkRR=>sbCG2R;
RRRRRRRRR#CDCR
RRRRRRRRRRVRss0NORR:=VOsN0R;
RRRRRRRRRsRRCRGbR=R:RbCG;R
RRRRRRRRRCRM8H
V;RRRRRRRRCCD#
RRRRRRRRsRRCRGbR=R:RbCG;R
RRRRRRRRRsNVsO:0R=FR50sEC#>R=R''j2R;
RRRRRRRRRssVNRO05NVsOF0HMH_I8-0E4FR8IFM0RNVsOF0HMH_I8-0E4N-5sHo_ME0'H-oE4R22:R=
RRRRRRRRRNRRsHo_M50RN_soH'M0EEHo-84RF0IMF2Rj;R
RRRRRRMRC8VRH;R
RRRRRRCRs#0kDRG5CbCFMMI0_HE802=R:Ro#HMR;
RRRRRCRRGMbFRR:=zQh1t7h RC5sG4b-2R;
RRRRRCRRGMbF5bCGFMMC0H_I8-0E4R2RRRRRRRRRR=R:R0MFRbCGFCM5GMbFC_M0I0H8E2-4;R
RRRRRRCRs#0kDRG5CbCFMMI0_HE80-84RF0IMF2RjRR:=z h)1emp V7_D0FN5bCGF;M2
RRRRRRRR#sCkRD05R-48MFI0-FRVOsN0MHF_8IH0RE2:z=Rh1) m pe7D_VF5N0sNVsO;02
RRRRCRRMH8RVR;
RCRRMH8RVR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-R8#0_oDFHPO_CFO0sFR0RFVDNR0
RMVkOF0HMFR0_FVDN50R
RRRRoNsRRRRRRRRRRRRRRRRRRRRR1:Raz7_pQmtB _eB)am;R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)Rqp:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820ER-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCVNbPsRR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RLHCoMR
RRVRHRoNs'MDCoR0E<RR40MEC
RRRRsRRCs0kMqRhw
u;RRRRCRM8H
V;RRRRVNbPs=R:R)zh p1me_ 7VNDF0s5No
2;RRRRskC0sVMRbsPN;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-RsbkbCF#:FROMsPC0N#RRHkVGRC80NFRRFVDNM0HoFRbH
M0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp k7_VCHG8R;R-k-RMo#HMRC8VCHG8FRbHRM0HkMb0R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)RqpR:RR=DRVF_N0CFGbM0CM_8IH0RE;RR--I0H8EVRFRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--I0H8EVRFRNVsOF0HMR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0M80RCsMFlHNDxRCRRRR:Apmm RqhR:RR=DRVF_N08FCMsDlNH2xCR-R-RCk#RCHCCGRC0#CMH#FM
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHND#CRNRsoRRR:#GVHC58RN'soEEHo+84RF0IMFsRNoF'DIR2;RR--1MHoCP8RCHs#FFMRVsRNoR
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RLHCoM-RR-kRVMHO0F0MRFD_VF
N0RRRRH5VRN'soDoCM0<ERRR420MEC
RRRRsRRCs0kMqRhw
u;RRRRCRM8H
V;RRRR#oNsRs5NoN'sM2oCRR:=#GVHC58RN2so;R
RRNR#s5oR#oNs'oEHE:2R=jR''R;
RsRRCD#k0=R:R_0FVNDF0NR5sRoRRRRRRRRRR>R=Rs#NoR,
RRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM0VF_D0FN;R

RMVkOF0HMFR0_FVDN50R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7V_#H8GC;RRRRR--#MHoCV8RH8GCRHbFMR0
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRRRR:V=RD0FN_bCGFMMC0H_I8;0ER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)RqpR:RR=DRVF_N0VOsN0MHF_8IH0RE;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0FRsk_M8#D0$CRRRRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHM
RRRRMOF#M0N0CR8MlFsNxDHCRRRRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--sMFk8oHMR0FbH
FMRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0MRH0CCosH_I8R0ERRRR:hRQa  t)=R:RoNs'oEHER;
RORRF0M#NRM0HVM_s0NOH_FMI0H8ERR:Q hatR ):N=RsDo'F
I;RRRRPHNsNCLDRCGs#0kDRRRRR#:RVCHG8HR5Mo0CCIs_HE80RI8FMR0FHVM_s0NOH_FMI0H8E
2;RRRRPHNsNCLDR#sCkRD0RRRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2
RRRRsPNHDNLCsRNoM_H0RRRRRR:zQh1t7h 50HMCsoC_8IH0-ERR_HMVOsN0MHF_8IH0-ERRR4
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR8RRF0IMF2Rj;-RR-HR#o8MCRsPC#MHFRRFVNksol0CM
RRRRsPNHDNLCsRNoRGRRRRRRRR:1hQt 57RHCM0o_CsI0H8ERR-HVM_s0NOH_FMI0H8EFR8IFM0R;j2
RRRRsPNHDNLCGRCbC,RGlb0bRR:1hQt 57RCFGbM0CM_8IH08ERF0IMF2Rj;R
RRNRPsLHNDCCRGMbFRRRRR:RRR1zhQ th7CR5GMbFC_M0I0H8ERR-4FR8IFM0R;j2
RRRRR--zHM#o8MCRsPC#MHFRRFVC3Gb
RRRRMOF#M0N0GRCb_FMLCN#RRR:1hQt 57RCFGbM0CM_8IH04E-RI8FMR0Fj:2R=R
RRRRRo_CMCFGbMN_L#CC5GMbFC_M0I0H8ER2;R-R-RbCGFMMC0VRFV0#C
RRRRsPNHDNLCsRVN,O0RNVsOl00bRR:zQh1t7h Rs5VNHO0FIM_HE80-84RF0IMF2RjR
:=RRRRRFR50sEC#>R=R''j2R;
RPRRNNsHLRDCsMFk8RR:Apmm Rqh:V=RNCD#;R
RLHCoMR
RRVRHRs5NoC'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMhuqw;R
RRMRC8VRH;R
RRsRGCD#k0=R:R_0FjN45sRo,'2X';R
RRsRNoRGRR=R:Rt1Qh5 70#F_DGP5skC#D202;R
RRVRHR#5Q_5XRN2so2ER0CRM
RRRRR#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRCHD#VNR5sRoG=2RjRC0EMR
RRRRRskC#D:0R=FR50sEC#>R=R''j2R;
RCRRD
#CRRRRRCRs#0kDRR:=5EF0CRs#='>Rj;'2RRRRRRRR-x-RCRsFFRk00RECskC#DR0
RRRRRRHVNGso5oNsGC'DVR02=4R''ER0CRMRR-RR-FR0#0#RE#CRHRoML
H0RRRRRRRRskC#D50RCFGbM0CM_8IH0RE2:'=R4R';RRRR-h-RC0oNHRPCMLklCRs
RRRRRNRRsRoGRRRRRRRRRRRRRRRRR:RR=NR-s;oGR-RR-NRv	HCR0FRb#HH0P
C3RRRRRDRC#RC
RRRRRsRRCD#k0CR5GMbFC_M0I0H8E:2R=jR''R;
RRRRR8CMR;HV
RRRRNRRsHo_M:0R=hRz1hQt 075Fj_G4a517m_pt_QBea Bm5)RNGso5oNs_0HM'MsNo2C22
2;RRRRR-R-RlBFbCk0Rb GFMMC0R
RRRRRCRGbRRRR:0=RFH_#o8MC5MVH8C_DVF0l#N05sHo_MR0,'24',GRCbC'DMEo02R;R-p-RF
o.RRRRRVRHRbCGRH+RMs_VNHO0FIM_HE80RC>RGMbF_#LNCER0CRMR-s-RCs0kMMRHVHHM0R$
RRRRRsRRCD#k0-R54FR8IFM0Rs-VNHO0FIM_HE802:RR=FR50sEC#>R=R''j2R;
RRRRRsRRCD#k0CR5GMbFC_M0I0H8E4R-RI8FMR0Fj:2R=FR50sEC#>R=R''42R;
RRRRRsRRCs0kMCRs#0kD;R
RRRRRCHD#V8R5CsMFlHNDxNCRMR8
RRRRRRRRRRRR5bCGRH+RMs_VNHO0FIM_HE80RR<=-#sCH5xCCFGbMN_L#RC,C'GbDoCM02E22ER0CRM
RRRRRCRRG:bR=sR-Cx#HCG5Cb_FMLCN#,GRCbC'DMEo02R;
RRRRR-RR-ER#HRV0LN$RRMOF#M0N0R
RRRRRRsRNoM_H0=R:RH#EVD0_CRV05oNs_0HM,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRs5NoM_H0H'Eo+ERR_0FHCM0o5CsCFGbMN_L#
C2RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR+MRH_NVsOF0HMH_I8R0E-2R42R;
RRRRRHRRVNR5sHo_ME0'HRoE>sRVNHO0FIM_HE802ER0CRM
RRRRRRRRRNVsO:0R=sRNoM_H0NR5sHo_ME0'H-oE4FR8IFM0Rs5NoM_H0H'EoVE-s0NOH_FMI0H8E;22
RRRRRRRRsRRF8kMRR:=OOEC	F_skRM85R
RRRRRRRRRRsRVN_O0HRMRR>R=RoNs_0HM5oNs_0HM'oEHEs-VNHO0FIM_HE802R,
RRRRRRRRR#RRHRoMRRRRR=RR>CRs#0kD5#sCk'D0EEHo2R,
RRRRRRRRRsRRCHlNMs8CR=RR>sRNoM_H0N55sHo_ME0'H-oEVOsN0MHF_8IH04E-2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2,RRRRRRRRRRRRsMFk80_#$RDC=s>RF8kM_$#0D;C2
RRRRRRRRHRRVsR5F8kM2ER0CRM
RRRRRRRRRVRRbF_skRM85NVsOH0_M>R=RoNs_0HMRs5NoM_H0H'Eo4E-RI8FM
0FRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR5RRN_soH'M0EEHo-NVsOF0HMH_I820E2R,
RRRRRRRRRRRRRRRRRRRRRbCGFHM_M=RR>GRCbR,
RRRRRRRRRRRRRRRRRRRRRNVsOF0_k=0R>sRVN,O0
RRRRRRRRRRRRRRRRRRRRCRRGMbF_0FkRR=>C0Gbl;b2
RRRRRRRRRRRRbCGRR:=C0Gbl
b;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RC
RRRRRRRRRNVsO50RVOsN0MHF_8IH04E-RI8FMR0FVOsN0MHF_8IH04E--s5NoM_H0H'Eo4E-2:2R=R
RRRRRRRRRRsRNoM_H0NR5sHo_ME0'H-oE4FR8IFM0R;j2
RRRRRRRR8CMR;HV
RRRRCRRD
#CRRRRRRRRN_soHRM0:#=RE0HV_VDC0NR5sHo_MR0,N_soH'M0EEHo-_0FHCM0o5CsC2Gb2R;
RRRRRCRRGRbRR:RR=GRCbRR+HVM_s0NOH_FMI0H8ER;
RRRRRHRRVNR5sHo_ME0'HRoE>sRVNHO0FIM_HE802ER0CRM
RRRRRRRRRNVsO:0R=sRNoM_H0NR5sHo_ME0'H-oE4FR8IFM0Rs5NoM_H0H'EoVE-s0NOH_FMI0H8E;22
RRRRRRRRsRRF8kMRR:=OOEC	F_skRM85R
RRRRRRRRRRsRVN_O0HRMRR>R=RNVsOj052R,
RRRRRRRRR#RRHRoMRRRRR=RR>CRs#0kD5#sCk'D0EEHo2R,
RRRRRRRRRsRRCHlNMs8CR=RR>sRNoM_H0N55sHo_ME0'H-oEVOsN0MHF_8IH04E-2R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRI8FMR0Fj
2,RRRRRRRRRRRRsMFk80_#$RDC=s>RF8kM_$#0D;C2
RRRRRRRRHRRVsR5F8kM2ER0CRM
RRRRRRRRRVRRbF_skRM85NVsOH0_M=RR>sRVN,O0
RRRRRRRRRRRRRRRRRRRRCRRGMbF_RHMRR=>C,Gb
RRRRRRRRRRRRRRRRRRRRVRRs0NO_0FkRR=>VOsN0b0l,R
RRRRRRRRRRRRRRRRRRRRRCFGbMk_F0>R=RbCG02lb;R
RRRRRRRRRRsRVNRO0:V=Rs0NO0;lb
RRRRRRRRRRRRbCGR:RR=GRCbb0l;R
RRRRRRRRRCRM8H
V;RRRRRRRRCCD#
RRRRRRRRVRRs0NORs5VNHO0FIM_HE80-84RF0IMFsRVNHO0FIM_HE80-54-N_soH'M0EEHo-242R
:=RRRRRRRRRRRRN_soHRM05oNs_0HM'oEHER-48MFI0jFR2R;
RRRRRCRRMH8RVR;
RRRRR8CMR;HV
RRRRCRRGMbFRR:=zQh1t7h RC5s#CHx5bCG-R4,CFGbM0CM_8IH02E2;R
RRRRRCFGbMG5CbCFMMI0_HE80-R42RRRRRRRRR:RR=FRM0GRCb5FMCFGbM0CM_8IH04E-2R;
RRRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:z=Rh1) m pe7D_VF5N0CFGbM
2;RRRRRCRs#0kDR45-RI8FMR0F-NVsOF0HMH_I820ERR:=z h)1emp V7_D0FN5NVsO;02
RRRR8CMR;HV
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F0MRFD_VF;N0
R
R-#-RH_xCsRC#VOkM0MHF#R
R-Q-RMo0CC0sRFDRVF
N0RkRVMHO0F0MRFD_VFRN05R
RRsRNoRRRRRRRRRRRRRRRR:RRRaQh )t ;R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR2R-s-RF8kMHRMoFHb0FRM
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _FVDN50R#CHx_#sC'VDC0FR8IFM0Rx#HCC_s#H'so2E0;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0ssMRCD#k0R;
RCRRD
#CRRRRRCRs#0kDRR:=0VF_D0FNRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=Rx#HCC_s#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>-x#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D;C2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-RNsCDFR0RFVDNR0
RMVkOF0HMFR0_FVDN50R
RRRRoNsRRRRRRRRRRRRRRRRRRR:)p q;R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-z-R#QCR R  CCG0M88CR
wuRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7D_VFRN05x#HCC_s#C'DV80RF0IMFHR#xsC_Cs#'H0oE2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMskC#D
0;RRRRCCD#
RRRRsRRCD#k0=R:R_0FVNDF0NR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRRRRRRRRRRRRRRRRR8RRCsMFlHNDxRCRR>R=RM8CFNslDCHx2R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0F0MRFD_VF;N0
R
R-k-RMo#HMRC80VFRD0FN
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _1zhQ th7R;
R#RRH_xCsRC#RRRRRRRRRRRR:hRz)m 1p7e _FVDN
0;RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC2RR--sMFk8oHMR0FbH
FMRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7D_VFRN05x#HCC_s#C'DV80RF0IMFHR#xsC_Cs#'H0oE2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMskC#D
0;RRRRCCD#
RRRRsRRCD#k0=R:R_0FVNDF0NR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$2DC;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_FVDN
0;
-RR-HR#o8MCRR0FVNDF0R
RVOkM0MHFR_0FVNDF0
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;R
RRHR#xsC_CR#RRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR2R-s-RF8kMH
MoRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7D_VFRN05x#HCC_s#C'DV80RF0IMFHR#xsC_Cs#'H0oE2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMskC#D
0;RRRRCCD#
RRRRsRRCD#k0=R:R_0FVNDF0NR5sRoRRRRRRRRRR>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F
I,RRRRRRRRRRRRRRRRRRRRRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$2DC;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_FVDN
0;
-RR-0R#8D_kFOoH_OPC0RFs0VFRD0FN
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRR:aR17p_zmBtQ_Be a;m)
RRRRx#HCC_s#RR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0#R5H_xCs'C#D0CVRI8FMR0F#CHx_#sC'osHE;02
LRRCMoH
RRRRRHV5#sCk'D0DoCM0<ERRR420MEC
RRRRsRRCs0kMCRs#0kD;R
RRDRC#RC
RRRRR#sCkRD0:0=RFD_VFRN05oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=->R#CHx_#sC'IDF2R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0F0MRFD_VF;N0
R
R-k-RMo#HMRC8VCHG8FRbHRM00VFRD0FN
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _HkVG;C8R-R-R#kMHCoM8HRVGRC8bMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HoR
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RkCCRHCCCRGM0C#MHF#R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0#R5H_xCs'C#D0CVRI8FMR0F#CHx_#sC'osHE;02
LRRCMoH
RRRRRHV5#sCk'D0DoCM0<ERRR420MEC
RRRRsRRCs0kMCRs#0kD;R
RRDRC#RC
RRRRR#sCkRD0:0=RFD_VFRN05oNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRRRRRNVsOF0HMH_I8R0E=->R#CHx_#sC'IDF,R
RRRRRRRRRRRRRRRRRRRRRRRRRsMFk80_#$RDCR=RR>FRsk_M8#D0$CR,
RRRRRRRRRRRRRRRRRRRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FVNDF0
;
R-R-Ro#HMRC8VCHG8FRbHRM00VFRD0FN
VRRk0MOHRFM0VF_D0FNRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _H#VG;C8
RRRRx#HCC_s#RRRRRRRRRRRRRR:z h)1emp V7_D0FN;R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MRo
RORRF0M#NRM08FCMsDlNHRxC:mRAmqp hRRRRR:=VNDF0C_8MlFsNxDHCR2R-s-RF8kMHRMoFHb0FRM
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _FVDN50R#CHx_#sC'VDC0FR8IFM0Rx#HCC_s#H'so2E0;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0ssMRCD#k0R;
RCRRD
#CRRRRRCRs#0kDRR:=0VF_D0FNRs5NoRRRRRRRRRRRRR=>N,so
RRRRRRRRRRRRRRRRRRRRRRRRCRRGMbFC_M0I0H8E>R=Rx#HCC_s#H'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>-x#HCC_s#F'DIR,
RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRCR8MlFsNxDHCRRRRR=>8FCMsDlNH2xC;R
RRRRRskC0ssMRCD#k0R;
RCRRMH8RVR;
R8CMRMVkOF0HMFR0_FVDN
0;
-RR-FR0_0HMCsoCRD5VF2N0
VRRk0MOHRFM0HF_Mo0CC5sR
RRRRoNsRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;RRR-V-RD0FNHRMobMFH0MRHb
k0RRRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs2FsR-R-RCOEOV	RFCsRsssF#R
RRCRs0MksRaQh )t 
HRR#R
RRNRPsLHNDPCRN8DHV:bRRDPNHV8_bN#00RC;R-R-RDeNHw8Ru0R#N
0CRRRRPHNsNCLDRNVsORRRRz:Rht1QhR 75s-NoF'DIFR8IFM0R;j2RRRRRRRRRR--wOsN0MHF
RRRRsPNHDNLCsRVN,O0RNVsO00_lRbRRz:Rht1QhR 75N4-sDo'F8IRF0IMF2Rj;RRRRRRRRR--wOsN0MHF
RRRRsPNHDNLCGRCbRFMRRR:1hQt 57RN'soEEHo-84RF0IMF2Rj;R
RRNRPsLHNDHCR#MHoR:RRR71a_mzpt;QBRRRRR-R-R0HMCNsMDCRPsF#HMVRFRo#HMR
RRNRPsLHNDsCRF8kMR:RRR71a_mzpt;QBRRRRR-R-RRH#sMFk8oHMRCMC8?C8
RRRRsPNHDNLCCRs#0kDRRR:Q hat; )
RRRRsPNHDNLCNRL#RCRRRR:Q hat; )RRRRRRRRRR--QCM0oRCsCFGbM0CM
RRRRsPNHDNLC0R#NHs08:GRR0HMCsoCRMsNoVCRs'NOEEHoRI8FMR0FjR;
RPRRNNsHLRDCskC8OeC8C:O0R8#0_FkDo;HO
LRRCMoH
RRRRDPNHb8VRR:=O#DN#RVb5oNs,EROC_O	CFsss
2;RRRRO#DN##ONCRR:OCN#RDPNHb8VR
H#RRRRRERICHMR#|GRRMMNRJ|Rk0HC_MMNRb|RFx#_CRsF|CRMoC_xs|FRR#bF_M8CFNslDRR|M_Co8FCMsDlNR
=>RRRRRRRRskC#D:0R=;RjRRRRRRRRRRRRRRRRRRRR-s-RCs0kM
RjRRRRRERICbMRFH#_M=VR>R
RRRRRRCRs#0kDRR:=Q hat' )EEHo;R
RRRRRIMECRoMC_VHMR
=>RRRRRRRRskC#D:0R=hRQa  t)F'DIR;
RRRRRCIEM0RFE#CsR
=>RRRRRRRRLNsC	k_MlsLCRR5
RRRRRRRRRoNsRRRRRRRRRR=>N,so
RRRRRRRRVRRbb0$RRRRR=RR>NRPDVH8bR,
RRRRRRRRRM8CFNslDCHxRR=>V#NDCR,
RRRRRRRRRNVsOR0RRRRRRR=>VOsN,R
RRRRRRRRRCFGbMRRRRRRR=C>RGMbF2R;
RRRRRVRRs0NORs5VN'O0EEHo2RRRRRRRRRRRRR:=';j'R-R-R8q8R0CGsLNRHV0RFjsR3OnRN
#CRRRRRRRRVOsN0VR5s0NO'oEHER-48MFI0jFR2=R:RNVsOR;
RRRRRHRR#MHoRRRRRRRRRRRRRRRRRRRRRRRRRR:=0GF_j54RNRso5oNs'oEHE;22
RRRRRRRR#LNCRRRRRRRRRRRRRRRRRRRRRRRR:RR=FR0_0HMCsoCRG5Cb2FMR4+R;R
RRRRRRVRHR#LNCRR<-04RE
CMRRRRRRRRRCRs#0kDRR:=jR;
RRRRRCRRDV#HR#LNC=R>RNVsOH'Eo0ERE
CMRRRRRRRRRCRs#0kDRR:=0HF_Mo0CC5sRVOsN0*2RR*.*5#LNCRR-VOsN'oEHE
2;RRRRRRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRR-W-RCCRMC08RFFRsk
M8RRRRRRRRRVRHR#LNCRR=-04RERCMRRRRRRRRRRRR-0-RsRNbVRFsjR3nOCN#3R
RRRRRRRRRRCRs#0kDRR:=jR;
RRRRRRRRR#CDCR
RRRRRRRRRR-RR-I)CsCH0RC0ERDVFDHFIMDoRHRMCFOVRFR8C0lFRNR	C#0$MEHC#xDNLCNR5P8FHRsCsF#sRNM$HoR
RRRRRRRRRR-RR-FRMMF-OMN#0MH0RMG8CRRHM#ODHCCRLO#NkCVRFRs"VNEO'H-oELCN#"RRRRZheRm.-Oj0-gR
RRRRRRRRRR-RR-#sCkRD0:0=RFM_H0CCosVR5s0NORs5VNEO'HRoE8MFI0VFRs'NOEEHo-#LNC;22
RRRRRRRRRRRRRRRVOsN0l_0b=R:RNVsO#0Rs5DRVOsN'oEHERR-LCN#2R;
RRRRRRRRRRRRRCRs#0kDRR:=0HF_Mo0CCVs5s0NO_b0l2R;
RRRRRRRRRRRR-C-RMF8RVCRsI0sHCR
RRRRRRRRRCRM8H
V;RRRRRRRRR-R-RksFMM8HoFRskM0HCR
RRRRRRRRROCN#RksFM#8_0C$DR
H#RRRRRRRRRRRRIMECRksFMM8_CCNs#=0R>R
RRRRRRRRRRRRRHVVRs'NOEEHoRL-RNR#C>RR40MEC
RRRRRRRRRRRRRRRR)--CHIs00CREVCRFFDDIoHMRDdRH#MCRRFVOCF8RR0FlCN	RM#$0#ECHLxND5CRNHPF8sRCsRFs#HN$MRo
RRRRRRRRRRRRR-RR-FRMMF-OMN#0MH0RMG8CRRHM#ODHCCRLO#NkCVRFRs"FRs5VNRO05NVsOH'Eo-ERR#LNCRR-.FR8IFM0R2j2"RRRRZheRm4-Oj0-gR
RRRRRRRRRRRRRR-R-sMFk8=R:RNVsO50RVOsN'oEHERR-LCN#R4-R2MRN8R
RRRRRRRRRRRRRR-R-RRRRRRRRRs5VNRO05NVsOH'Eo-ERR#LNCR2
RRRRRRRRRRRRR-RR-RRRRRRRRFRRsFR5sVR5s0NORs5VNEO'HRoE-NRL#-CRR8.RF0IMF2Rj2;22
RRRRRRRRRRRRRRRRN#0s80HG=R:RNVsOH'Eo-ERR#LNCRR-.R;
RRRRRRRRRRRRRsRRCO8kCC8eO:0R=jR''R;
RRRRRRRRRRRRRVRRFQsRRRHMVOsN0Q']t8]RF0IMFRRjDbFF
RRRRRRRRRRRRRRRRRRRRRHVQ=R<RN#0s80HGER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRskC8OeC8CRO0:s=RCO8kCC8eOF0RssRVN5O0Q
2;RRRRRRRRRRRRRRRRRRRRCRM8HRV;
RRRRRRRRRRRRRRRR8CMRFDFbR;
RRRRRSRSSRR
RRRRRRRRRRRRRsRRF8kMRR:=VOsN0VR5s'NOEEHoRL-RNR#C-2R4R8NM
RRRRRRRRRRRRRRRRRRRRRRRRVR5s0NORs5VNEO'HRoE-NRL#RC2FssRCO8kCC8eO;02
RRRRRRRRRRRRRRRRR--CRM8FsVRCHIs0RC
RRRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRRFRskRM8:V=Rs0NORs5VNEO'HRoE-NRL#-CRRR42N
M8RRRRRRRRRRRRRRRRRRRRRRRRRNVsO50RVOsN'oEHERR-LCN#2R;
RRRRRRRRRRRRR8CMR;HV
RRRRRRRRRRRRCIEMFRsk_M8HRMV=R>
RRRRRRRRRRRRRksFM:8R=sRVN5O0VOsN'oEHERR-LCN#R4-R2MRN8FRM0#RHH;oM
RRRRRRRRRRRRCIEMFRsk_M8MHCoM=VR>R
RRRRRRRRRRRRRsMFk8=R:RNVsOV05s'NOEEHoRL-RNR#C-2R4R8NMRHH#o
M;RRRRRRRRRRRRIMECREF0CRs#=R>
RRRRRRRRRRRRRksFM:8R=jR''R;
RRRRRRRRR8CMR#ONCR;
RRRRRRRRRRHVsMFk8RR='R4'0MEC
RRRRRRRRRRRR#sCkRD0:s=RCD#k0RR+4R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
RRRRRRRRRHVHo#HMRR='R4'0MEC
RRRRRRRRsRRCD#k0=R:Rs-RCD#k0R;
RRRRRCRRMH8RVR;
RCRRMO8RNR#CO#DN##ONCR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FHCM0o;Cs
R
R-0-RFM_k#MHoC58RVNDF0R2
RMVkOF0HMFR0_#kMHCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRR:RRRahqzp)q;RRRR-R-RMDCoR0EFFVRkk0b0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF2-RR-EROCRO	VRFsCFsssR#
RsRRCs0kMhRz)m 1p7e _1zhQ th7R
RHR#
RPRRNNsHLRDCPHND8RVb:NRPD_H8V0b#N;0CR-RR-NReDRH8w#uR0CN0
RRRRsPNHDNLCsRVNRORRRR:z h)1emp z7_ht1QhR 75x#HCR-48MFI0jFR2R;R-w-Rs0NOH
FMRRRRPHNsNCLDRo#HMRRRR1:Raz7_pQmtBR;RRRRR-M-RFk0R#
C8RCRLo
HMRRRRPHND8RVb:O=RD#N#V5bRN,soRCOEOC	_sssF2R;
RORRD#N#OCN#RO:RNR#CPHND8RVbHR#
RRRRRCIEM#RHGRR|MRNM|kRJH_C0MRNM=R>
RRRRRVRRsRNO:5=RFC0Es=#R>XR''
2;RRRRRERICbMRFx#_CRsF|CRMoM_HVRR|M_CoxFCsRM|RCMo_FNslDRR|b_F#8FCMsDlNRM|RC8o_CsMFlRND=R>
RRRRRVRRsRNO:5=RFC0Es=#R>jR''R2;RRRRR-RR-CRs0MksRRj
RRRRRCIEMFRb#M_HV>R=
RRRRRRRRNVsO=R:R05FE#CsRR=>'24';R
RRRRRIMECREF0CRs#=R>
RRRRRVRRD0FN__0FkHM#o8MCRR5
RRRRRRRRRoNsRRRRRRRRRR=>N,so
RRRRRRRRVRRsRNORRRRR=RR>sRVN
O,RRRRRRRRRHR#oRMRRRRRR>R=Ro#HMR,
RRRRRRRRRM8CFNslDCHxRR=>V#NDCR,
RRRRRRRRRNLH#RRRRRRRRR=>jR,
RRRRRRRRRksFM#8_0C$DRR=>sMFk80_#$2DC;R
RRMRC8NRO#OCRD#N#OCN#;R
RRCRs0MksRs5VN;O2
CRRMV8Rk0MOHRFM0kF_Mo#HM;C8
R
R-0-RFH_#o8MCRD5VF2N0
VRRk0MOHRFM0#F_HCoM8
R5RRRRNRsoRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRFROMN#0M#0RHRxCRRRRR:RRRahqzp)q;RRRR-R-RMDCoR0EFFVRkk0b0R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF2-RR-EROCRO	VRFsCFsssR#
RsRRCs0kMhRz)m 1p7e _t1Qh
 7R#RH
RRRRsPNHDNLCHR#oRMRRRR:1_a7ztpmQRB;RRRRRR--0CskRRHVMNCo0CHP
RRRRsPNHDNLCNRPDVH8bRR:PHND8b_V#00NCR;RRR--eHND8uRwRN#00RC
RPRRNNsHLRDCVOsNRRRR:hRz)m 1p7e _1zhQ th7#R5H-xC4FR8IFM0R;j2R-R-RNwsOF0HMR
RRNRPsLHNDsCRCD#k0:RRR)zh p1me_ 71hQt 57R#CHx-84RF0IMF2Rj;R
RLHCoMR
RRNRPDVH8b=R:RNOD#b#VRs5NoO,RE	CO_sCsF;s2
RRRRNOD#N#O#:CRR#ONCNRPDVH8b#RH
RRRRIRRERCMHR#G|NRMMRR|JCkH0N_MM>R=
RRRRRRRR#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRRERICbMRFx#_CRsF|CRMoC_xs|FRR#bF_M8CFNslDRR|M_Co8FCMsDlNR
=>RRRRRRRRskC#D:0R=FR50sEC#>R=R''j2R;RRRRR-s-RCs0kM
RjRRRRRERICbMRFH#_M=VR>R
RRRRRRCRs#0kDRRRRRRRRRRRRR:RR=FR50sEC#>R=R''42R;
RRRRRsRRCD#k0sR5CD#k0H'EoRE2:'=Rj
';RRRRRERICMMRCHo_M=VR>R
RRRRRRCRs#0kDRRRRRRRRRRRRR:RR=FR50sEC#>R=R''j2R;
RRRRRsRRCD#k0sR5CD#k0H'EoRE2:'=R4
';RRRRRERICFMR0sEC#>R=
RRRRRRRRFVDN00_FM_k#MHoC58R
RRRRRRRRNRRsRoRRRRRR=RR>sRNoR,
RRRRRRRRRo#HMRRRRRRRRR=>#MHo,R
RRRRRRRRRVOsNRRRRRRRR=V>Rs,NO
RRRRRRRR8RRCsMFlHNDx=CR>NRVD,#C
RRRRRRRRLRRHRN#RRRRR=RR>,Rj
RRRRRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$C
2;RRRRRRRRskC#D50R#CHx-R42RRRRRRRRRR:=';j'
RRRRRRRR#sCkRD05x#HCR-.8MFI0jFR2=R:R)zh p1me_ 71hQt V75sRNO5x#HCR-.8MFI0jFR2
2;RRRRRRRRH#VRHRoM=4R''ER0CRM
RRRRRRRRRR--ANCOkR#C0RECl0F#RoMCNP0HCHR#o8MCRlMkLRCsH4#RR#DC#ER0N0MRElCRF
#0RRRRRRRRR-R-R#bFHP0HCHR#o8MCRlMkL,CsRRICM8CCRH0E#FRO8
C3RRRRRRRRRVRHRNVsOs5VNEO'H2oER'=R40'RERCMRRRRR-R-R0sCkRsMl0F#RoMCNP0HCkRMlsLC
RRRRRRRRRRRR#sCkRD0RRRRRRRRRRRRR=R:R05FE#CsRR=>'2j';R
RRRRRRRRRRCRs#0kDRC5s#0kD'oEHE:2R=4R''R;
RRRRRRRRR#CDCR
RRRRRRRRRRCRs#0kDRR:=-#sCk;D0
RRRRRRRRCRRMH8RVR;
RRRRRCRRD
#CRRRRRRRRRVRHRNVsOs5VNEO'H2oER'=R40'RERCMRRRRR-R-R0sCkRsMl0F#R#bFHP0HCkRMlsLC
RRRRRRRRRRRR#sCkRD0RRRRRRRRRRRRR=R:R05FE#CsRR=>'24';R
RRRRRRRRRRCRs#0kDRC5s#0kD'oEHE:2R=jR''R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
RRRR8CMR#ONCDRONO##N;#C
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F0MRFH_#o8MC;R

RR--bbksF:#CRMBFP0Cs#RRNVNDF0FR0RHkVG
C8RkRVMHO0F0MRFV_kH8GCRR5
RNRRsRoRRRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRRRRRRRRR-R-RRVbHkMb0R
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )R-R-R0HMCsoCRsbN0R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hat; )R-R-RNVsOF0HMNRbsR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0DRC;RR--#kN0sCN0
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR;R-s-RF8kMH
MoRRRRO#FM00NMRCOEOC	_sssFRRRR:mRAmqp hRRRRRRRRRRRRRRRRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxCR:RRRmAmph qRRRRRRRRRRRRRRRRR:RR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMz h)1emp k7_VCHG8R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRaQh )t RR:=-MlHCs5NoF'DIN,RsDo'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERR:Q hatR ):N=RsEo'H;oER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0M#0RHRxCRRRRRRRRRRR:Q hatR ):D=RC_V0HCM8GRR-sEHo0M_H8RCG+;RcR-R-R#kMHCoM8HR#xRC
RPRRNNsHLRDCCFGbMN_L#RCRR:RRRaQh )t ;-RR-GRCbCFMMF0RVCV#0R
RRNRPsLHNDPCRN8DHVRbRRRRRRRR:PHND8b_V#00NCR;RRRRRRRRRRRRRRR--eHND8uRwRN#00RC
RPRRNNsHLRDCCRGbRRRRRRRRR:RRRaQh )t ;-RR-GR bCFMMR0
RPRRNNsHLRDCCFGbMRRRRRRRR:RRR1zhQ th7CR5GMbFC_M0I0H8ER-48MFI0jFR2R;R-e-RCFO0sCHx8GRCbCFMMR0
R-RR-NRA#0CRFHR8PCH8RNVsOF0HM$RL
RRRRsPNHDNLCsRVNRORRRRRRRRRRz:Rht1QhR 75x#HCR-48MFI0jFR2=R:R05FE#CsRR=>'2j';-RR-sRwNHO0FRM
RPRRNNsHLRDCVOsN_H#EVR0RR:RRR1zhQ th7#R5H-xC4FR8IFM0R;j2R-R-RNwsOF0HMER#HCV08R
RRNRPsLHND#CRE0HVRRRRRRRRRRR:Q hat; )
RRRRsPNHDNLCCRs#0kD_oLHRRRRRz:Rh1) m pe7V_kH8GCRC5DVH0_MG8CRI8FMR0FsEHo0M_H8-CGd
2;RRRRPHNsNCLDR#sCkRD0RRRRRRRR:hRz)m 1p7e _HkVGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMC;G2R-R-R#sCk
D0RCRLoRHMRR--VOkM0MHFR_0FkGVHCR8
RPRRN8DHV:bR=DRONV##bNR5sRo,OOEC	s_Cs2Fs;R
RRDRONO##NR#C:NRO#PCRN8DHVHbR#R
RRRRRIMECRGH#RM|RN|MRRHJkCM0_N=MR>R
RRRRRRsRVN:OR=FR50sEC#>R=R''X2R;
RRRRRCIEMFRb#C_xs|FRRoMC_VHMRM|RCxo_CRsF|CRMoF_MsDlNRM|RC8o_CsMFlRND=R>
RRRRRVRRsRNO:5=RFC0Es=#R>jR''R2;RRRRR-RR-CRs0MksRRj
RRRRRCIEMFRb#M_HV>R=
RRRRRRRRNVsO=R:R05FE#CsRR=>'24';RRRRRRRRR--NNDI$##RNs0kN
0CRRRRRERICFMR0sEC#>R=
RRRRRRRRbCGFLM_NR#C:.=R*C*5GMbFC_M0I0H8E2-4R;-4RRRRRRRRRRRR-C-RGMbFCRM0F#VVCR0
RRRRR-RR-HRwoCksR0FkRC0ERNVsOF0HMR
RRRRRRVRHRN5PDVH8bRR=b_F#8FCMsDlN2MRN8CR8MlFsNxDHCER0CRM
RRRRRRRRRbCGRRRRRRRRRRRRR=R:RG-Cb_FMLCN#R;+4
RRRRRRRRVRRsRNO5NVsOH'EoRE2:'=RjR';RRRRRR--)FClP0CRE"CR4"3j3R
RRRRRRDRC#RC
RRRRRRRRRR--CFGbM0CMRR/=',j'RsMFlRNDVNDF0oHMRHbFMR0
RRRRRRRRRbCGFRMRRRRRRRRRRRRRRRRRRR:=zQh1t7h 5oNsRG5CbCFMMI0_HE80-84RF0IMF2Rj2R;
RRRRRRRRRbCGFCM5GMbFC_M0I0H8E2-4RR:=MRF0CFGbMG5CbCFMMI0_HE80-;42
RRRRRRRRCRRGRbRRRRRRRRRRRRRRRRRR:RR=FR0_0HMCsoCRQ51t7h 5bCGF2M2R;+4
RRRRRRRRVRRsRNO5NVsOH'EoRE2RRRRR:RR=4R''R;RRR--qR880REC"j43"R3
RRRRRCRRMH8RVR;
RRRRR#RRE0HVRR:=5NVsOH'Eo-ERR+dRRosHEH0_MG8C2RR-C;Gb
RRRRRRRRRHVVOsN0MHF_8IH0>ERRNVsOH'Eo0ERERCMRR--BRNMF$MDRCk#Rx#HCR-.L#H0
RRRRRRRRVRRsRNO5NVsOH'Eo4E-RI8FMR0Fj:2R=hRz1hQt 57R0#F_D5PRN5so-84RF0IMFR
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRs-VNEO'H2oE2
2;RRRRRRRRCCD#RRRRRRRRRRRRRRRRRRRRRRRRRRRR-O-RNkMR#NCRDLDRH
0#RRRRRRRRRsRVN5ORVOsN'oEHER-48MFI0VFRs'NOEEHo-NVsOF0HMH_I820ER
:=RRRRRRRRRRRRzQh1t7h RF50_P#DRs5No45-RI8FMR0F-NVsOF0HMH_I820E2
2;RRRRRRRRCRM8H
V;RRRRRRRRVOsN_H#EV:0R=sRVN#ORs#DRE0HV;R
RRRRRRVRHRH#EV<0RR0jRERCMRRRRRRRRRRRRR-R-RCmPsFVDIR
RRRRRRRRRVOsNRR:=5EF0CRs#='>R4;'2
RRRRRRRR#CDCR
RRRRRRRRRVOsNRR:=VOsN_H#EV
0;RRRRRRRRCRM8H
V;RRRRCRM8OCN#RNOD#N#O#
C;RRRRskC#DL0_H:oR=FR0_HkVGRC85R
RRRRRNRsoRRRRRRRR=1>Raz7_pQmtB _eB)am5NVsO
2,RRRRRCRDVH0_MG8CR>R=RVDC0M_H8,CG
RRRRsRRH0oE_8HMC=GR>sR5H0oE_8HMCdG-2
2;RRRRskC#D:0R=CRs#CHxRs5NoRRRRRRRRRRRRR=>skC#DL0_H
o,RRRRRRRRRRRRRRRRRRRRRCRDVH0_MG8CRRRRRR=>D0CV_8HMC
G,RRRRRRRRRRRRRRRRRRRRRHRso_E0HCM8GRRRRR=>sEHo0M_H8,CG
RRRRRRRRRRRRRRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRRRRRRFsPCVIDF_$#0D=CR>PRFCDsVF#I_0C$D2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0FkGVHC
8;
-RR-kRbs#bFCB:RFCMPsR0#NDRVFRN00#FRVCHG8R
RVOkM0MHFR_0F#GVHC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RRVbHkMb0R
RRFROMN#0MD0RC_V0HCM8GRRRRRR:Q hat; )R-R-R0HMCsoCRsbN0R
RRFROMN#0Ms0RH0oE_8HMCRGRRRR:Q hat; )R-R-RNVsOF0HMNRbsR0
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0DRC;RR--#kN0sCN0
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR;R-s-RF8kMH
MoRRRRO#FM00NMRCOEOC	_sssFRRRR:mRAmqp hRRRRRRRRRRRRRRRRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxCR:RRRmAmph qRRRRRRRRRRRRRRRRR:RR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RORRF0M#NRM0VOsN0MHF_8IH0:ERRaQh )t RR:=-MlHCs5NoF'DIN,RsDo'F;I2R-R-RMDCoR0EFwVRukRF00bkRNVsOF0HMR
RRFROMN#0MC0RGMbFC_M0I0H8ERR:Q hatR ):N=RsEo'H;oER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRFROMN#0M#0RHRxCRRRRRRRRRRR:Q hatR ):D=RC_V0HCM8GRR-sEHo0M_H8RCG+;RcR-R-R#kMHCoM8HR#xRC
RPRRNNsHLRDCCFGbMN_L#RCRR:RRRaQh )t ;-RR-GRCbCFMMF0RVCV#0R
RRNRPsLHNDPCRN8DHVRbRRRRRRRR:PHND8b_V#00NCR;RR-RR-NReDRH8w#uR0CN0
RRRRsPNHDNLCGRCbRRRRRRRRRRRRQ:Rhta  R);RR-- FGbM0CM
RRRRsPNHDNLCHR#oRMRRRRRRRRRRA:Rm mpqRh;RR--0CskRRHVMNCo0CHP
RRRRsPNHDNLCGRCbRFMRRRRRRRRRz:Rht1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2R-R-ROeC0HFsxRC8CFGbM0CM
RRRRR--ACN#RR0F8HHP8VCRs0NOHRFMLR$
RPRRNNsHLRDCVOsNRRRRRRRRR:RRR1zhQ th7#R5H-xC.FR8IFM0RRj2:5=RFC0Es=#R>jR''R2;RR--wOsN0MHF
RRRRsPNHDNLCsRVN#O_E0HVRRRRRz:Rht1QhR 75x#HCR-.8MFI0jFR2R;R-w-Rs0NOHRFM#VEH0
C8RRRRPHNsNCLDRH#EVR0RRRRRRRRR:hRQa  t)R;
RPRRNNsHLRDCso#HMRC8RRRRR:RRRt1QhR 75x#HCR-48MFI0jFR2R;R-#-RHCoM8CRPsF#HMVRFR#sCk
D0RRRRPHNsNCLDR#sCk_D0LRHoRRRR:hRz)m 1p7e _H#VGRC85VDC0M_H8RCG8MFI0sFRH0oE_8HMCdG-2R;
RPRRNNsHLRDCskC#DR0RRRRRR:RRR)zh p1me_ 7#GVHC58RD0CV_8HMC8GRF0IMFHRso_E0HCM8GR2
RRRRRR:=5EF0CRs#='>Rj;'2R-R-R#sCk
D0RCRLoRHMRR--VOkM0MHFR_0F#GVHCR8
RPRRN8DHV:bR=DRONV##bNR5sRo,OOEC	s_Cs2Fs;R
RRDRONO##NR#C:NRO#PCRN8DHVHbR#R
RRRRRIMECRGH#RM|RN|MRRHJkCM0_N=MR>R
RRRRRRCRs#0kDRR:=5EF0CRs#='>RX;'2
RRRRIRRERCMb_F#xFCsRM|RCxo_CRsF=R>
RRRRRsRRCD#k0=R:R05FE#CsRR=>'2j';RRRR-RR-CRs0MksRRj
RRRRRCIEMCRMoM_HV>R=
RRRRRRRR#sCkRD05VDC0M_H82CGRR:=';4'RRRRRR--skC0s#MRlDNDCR#0MNCo0CHPRlMkL
CsRRRRRERICbMRFH#_M=VR>R
RRRRRRCRs#0kDRRRRRRRRRRRRR=R:R05FE#CsRR=>'24';-RR-CRs0MksRsDNo0C#RlMkL
CsRRRRRRRRskC#D50RD0CV_8HMCRG2:'=Rj
';RRRRRERICFMR0sEC#>R=
RRRRRRRRbCGFLM_NR#C:.=R*C*5GMbFC_M0I0H8E2-4R;-4R-R-RbCGFMMC0VRFV0#C
RRRRRRRRRHVN5soCFGbM0CM_8IH0RE2=jR''ER0CRM
RRRRRRRRRo#HM=R:RDVN#
C;RRRRRRRRCCD#
RRRRRRRR#RRHRoM:0=Rs;kC
RRRRRRRR8CMR;HV
RRRRRRRRR--wkHosFCRk00REVCRs0NOH
FMRRRRRRRRH5VRPHND8RVb=FRb#C_8MlFsNFDRsNRPDVH8bRR=M_Co8FCMsDlN2R
RRRRRRRRRNRM88FCMsDlNHRxC0MEC
RRRRRRRRCRRGRbRRRRRRRRRRRRR:-=RCFGbMN_L#+CR4R;
RRRRRRRRRNVsOVR5s'NOEEHo2=R:R''j;RRRR-RR-8Rq8ER0C4R"33j"
RRRRRRRR#CDCR
RRRRRRRRR-C-RGMbFCRM0/'=RjR',MlFsNVDRD0FNHRMobMFH0R
RRRRRRRRRCFGbMRRRRRRRRRRRRRRRRRRR:z=Rht1Qh5 7NRso5bCGFMMC0H_I8-0E4FR8IFM0R2j2;R
RRRRRRRRRCFGbMG5CbCFMMI0_HE80-R42:M=RFC0RGMbF5bCGFMMC0H_I8-0E4
2;RRRRRRRRRGRCbRRRRRRRRRRRRRRRRRRRR=R:R_0FHCM0oRCs5t1Qh5 7CFGbMR22+
4;RRRRRRRRRsRVN5ORVOsN'oEHER2RRRRRR=R:R''4;RRRRRRRRR--qR880REC"j43"R3
RRRRRCRRMH8RVR;
RRRRR#RRE0HVRR:=5NVsOH'Eo-ERR+dRRosHEH0_MG8C2RR-C;Gb
RRRRRRRRRHVVOsN0MHF_8IH0>ERRNVsOH'Eo0ERERCMRRRRR-R-RMBNRDFM$#RkCHR#x.C-R0LH#R
RRRRRRRRRVOsNRs5VNEO'H-oE4FR8IFM0RRj2:z=Rht1QhR 75_0F#RDP5oNs5R-48MFI0RF
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRVR-s'NOEEHo2;22
RRRRRRRR#CDCRRRRRRRRRRRRRRRRRRRRRRRRRRRRR--ORNMkR#CNRDDL#H0
RRRRRRRRVRRsRNO5NVsOH'Eo4E-RI8FMR0FVOsN'oEHEs-VNHO0FIM_HE802=R:
RRRRRRRRRRRR1zhQ th70R5FD_#PNR5s-o54FR8IFM0Rs-VNHO0FIM_HE802;22
RRRRRRRR8CMR;HV
RRRRRRRRNVsOE_#HRV0:V=RsRNO#RsD#VEH0R;
RRRRRHRRVER#HRV0<RRj0MECRRRRRRRRRRRRR-RR-PRmCDsVFRI
RRRRRRRRRNVsO=R:R05FE#CsRR=>'24';R
RRRRRRDRC#RC
RRRRRRRRRNVsO=R:RNVsOE_#H;V0
RRRRRRRR8CMR;HV
RRRRRRRRRHVMRF0#MHoRC0EMR
RRRRRRRRRso#HMRC8:1=RQ th7j5""RR&VOsN2R;
RRRRRCRRD
#CRRRRRRRRR#RsHCoM8=R:R1-5Q th7j5""RR&VOsN2
2;RRRRRRRRCRM8H
V;RRRRRRRRskC#DL0_H:oR=FR0_H#VGRC85R
RRRRRRRRRNRsoRRRRRRRR=1>Rap7_mBtQ_Be a5m)so#HM2C8,R
RRRRRRRRRD0CV_8HMCRGR=D>RC_V0HCM8GR,
RRRRRRRRRosHEH0_MG8CRR=>5osHEH0_MG8C-2d2;R
RRRRRRCRs#0kDRR:=sHC#x5CRNRsoRRRRRRRRR=RR>CRs#0kD_oLH,R
RRRRRRRRRRRRRRRRRRRRRRRRRD0CV_8HMCRGRR=RR>CRDVH0_MG8C,R
RRRRRRRRRRRRRRRRRRRRRRRRRsEHo0M_H8RCGR=RR>HRso_E0HCM8GR,
RRRRRRRRRRRRRRRRRRRRRRRRRksFM#8_0C$DRRRR=s>RF8kM_$#0D
C,RRRRRRRRRRRRRRRRRRRRRRRRRPRFCDsVF#I_0C$DRR=>FsPCVIDF_$#0D;C2
RRRR8CMR#ONCDRONO##N;#C
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F0MRFV_#H8GC;R

RR--#CHx_#sCRsPC#MHF#R
R-V-RD0FNRR0FkHM#o8MC
VRRk0MOHRFM0kF_Mo#HMRC85R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7h_z1hQt 
7;RRRRO#FM00NMRksFM#8_0C$DRs:RF8kM_b0$C=R:RFVDNs0_F8kM_$#0DRC;RR--sMFk8oHMR0FbH
FMRRRRO#FM00NMRCOEOC	_sssFRA:Rm mpqRhRR=R:RFVDNO0_E	CO_sCsFRs2RR--OOEC	FRVssRCs#Fs
RRRR0sCkRsMz h)1emp z7_ht1Qh
 7R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7h_z1hQt 57R#CHx_#sC'MsNo;C2
LRRCMoH
RRRRRHV5Z1Q  _)1C'DMEo0Rj=R2ER0CRM
RRRRR0sCkRsMskC#D
0;RRRRCCD#
RRRRsRRCD#k0=R:R_0FkHM#o8MCRR5
RRRRRNRRsRoRRRRRR=RR>sRNoR,
RRRRR#RRHRxCRRRRR=RR>HR#xsC_CD#'C0MoER,
RRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$CR,
RRRRRORRE	CO_sCsF=sR>EROC_O	CFsss
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0kF_Mo#HM;C8
R
R-V-RD0FNRR0F#MHoCR8
RMVkOF0HMFR0_o#HMRC85R
RRsRNoRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;R-V-RD0FNHRMobMFH0MRHb
k0RRRR#CHx_#sCRRRRRRRRRRRRRz:Rh1) m pe7Q_1t7h ;R
RRFROMN#0Ms0RF8kM_$#0D:CRRksFM08_$RbC:V=RD0FN_ksFM#8_0C$D;-RR-FRskHM8MFoRbF0HMR
RRFROMN#0MO0RE	CO_sCsF:sRRmAmph qRRRR:V=RD0FN_COEOC	_sssF2-RR-EROCRO	VRFsCFsssR#
RsRRCs0kMhRz)m 1p7e _t1Qh
 7R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7Q_1t7h RH5#xsC_Cs#'NCMo2R;
RoLCHRM
RHRRV1R5Q_Z )' 1DoCM0=ERRRj20MEC
RRRRsRRCs0kMCRs#0kD;R
RRDRC#RC
RRRRR#sCkRD0:0=RFH_#o8MCRR5
RRRRRNRRsRoRRRRRR=RR>sRNoR,
RRRRR#RRHRxCRRRRR=RR>HR#xsC_CD#'C0MoER,
RRRRRsRRF8kM_$#0D=CR>FRsk_M8#D0$CR,
RRRRRORRE	CO_sCsF=sR>EROC_O	CFsss
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_HCoM8
;
R-R-RsbkbCF#:FRBMsPC0N#RRFVDN00RFMRk#MHoCV8RH8GCRHbFMR0
RMVkOF0HMFR0_HkVGRC85R
RRsRNoRRRRRRRRRRRRRRRRRRRRRR:z h)1emp V7_D0FN;-RR-bRVRbHMkR0
R#RRH_xCsRC#RRRRRRRRRRRRR:RRR)zh p1me_ 7kGVHC
8;RRRRO#FM00NMRCFPsFVDI0_#$RDC:HRVG_C8FsPCVIDF_$#0D0C_$RbC:V=RH8GC_CFPsFVDI0_#$;DCR-R-R0#Nk0sNCR
RRFROMN#0Ms0RF8kM_$#0DRCRRRR:VCHG8F_sk_M8#D0$C$_0bRCRR=R:RGVHCs8_F8kM_$#0DRC;RR--sMFk8oHM
RRRRMOF#M0N0EROC_O	CFsssRRRRA:Rm mpqRhRRRRRRRRRRRRRRRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRRRR:mRAmqp hRRRRRRRRRRRRRRRRRRR:V=RD0FN_M8CFNslDCHx2R
RRCRs0MksR)zh p1me_ 7kGVHCR8
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _HkVGRC85x#HCC_s#C'DV80RF0IMFHR#xsC_Cs#'H0oE2R;
RoLCHRM
RHRRVsR5CD#k0C'DMEo0R4<R2ER0CRM
RRRRR0sCkRsMskC#D
0;RRRRCCD#
RRRRsRRCD#k0=R:R_0FkGVHC58R
RRRRRRRRoNsRRRRRRRRRRRR=N>Rs
o,RRRRRRRRD0CV_8HMCRGRR=RR>HR#xsC_CE#'H,oE
RRRRRRRRosHEH0_MG8CRRRR=#>RH_xCs'C#D,FI
RRRRRRRRCFPsFVDI0_#$RDC=F>RPVCsD_FI#D0$CR,
RRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRREROC_O	CFsssRRRRR=>OOEC	s_Cs,Fs
RRRRRRRRM8CFNslDCHxRRRR=8>RCsMFlHNDx;C2
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FkGVHC
8;
-RR-DRVFRN00#FRHCoM8HRVGRC8bMFH0R
RVOkM0MHFR_0F#GVHC58R
RRRRoNsRRRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0R-R-RRVbHkMb0R
RRHR#xsC_CR#RRRRRRRRRRRRRRRR:z h)1emp #7_VCHG8R;
RORRF0M#NRM0FsPCVIDF_$#0D:CRRGVHCF8_PVCsD_FI#D0$C$_0b:CR=HRVG_C8FsPCVIDF_$#0DRC;RR--#kN0sCN0
RRRRMOF#M0N0FRsk_M8#D0$CRRRRV:RH8GC_ksFM#8_0C$D_b0$CRRRRR:=VCHG8F_sk_M8#D0$CR;R-s-RF8kMH
MoRRRRO#FM00NMRCOEOC	_sssFRRRR:mRAmqp hRRRRRRRRRRRRRRRRRRR:V=RD0FN_COEOC	_sssF;-RR-EROCRO	VRFsCFsssR#
RORRF0M#NRM08FCMsDlNHRxCR:RRRmAmph qRRRRRRRRRRRRRRRRR:RR=DRVF_N08FCMsDlNH2xC
RRRR0sCkRsMz h)1emp #7_VCHG8R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7#GVHC58R#CHx_#sC'VDC0FR8IFM0Rx#HCC_s#H'so2E0;R
RLHCoMR
RRVRHRC5s#0kD'MDCoR0E<2R4RC0EMR
RRRRRskC0ssMRCD#k0R;
RCRRD
#CRRRRRCRs#0kDRR:=0#F_VCHG8
R5RRRRRRRRNRsoRRRRRRRRR=RR>sRNoR,
RRRRRDRRC_V0HCM8GRRRR>R=Rx#HCC_s#H'Eo
E,RRRRRRRRsEHo0M_H8RCGR=RR>HR#xsC_CD#'F
I,RRRRRRRRFsPCVIDF_$#0D=CR>PRFCDsVF#I_0C$D,R
RRRRRRFRsk_M8#D0$CRRRRR=>sMFk80_#$,DC
RRRRRRRRCOEOC	_sssFRRRR=O>RE	CO_sCsF
s,RRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHC
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0#F_VCHG8
;
R-R-R_0FsDCNRD5VF2N0
-RR-$R0bNHODRD$MRF010$MEHC#xDNLCMRkD#C#RC0ERbHMkH0R#RRNO#FM00NM3R
RVOkM0MHFR_0FsDCNRR5
RNRRsRoRRRRRRRRRRRRRRRRR:hRz)m 1p7e _FVDNR0;RRRRR-RR-DRVFHN0MboRF0HMRbHMkR0
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsM)p q
HRR#R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:Q hatR ):-=RlCHM5oNs'IDF,sRNoF'DIR2;RR--DoCM0FERVuRwR0FkbRk0VOsN0MHF
RRRRMOF#M0N0GRCbCFMMI0_HE80RQ:Rhta  :)R=sRNoH'EoRE;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRsPNHDNLCHR#oRMRRRRRRRRRR):R ;qpRRRRRR--1MHo,RR+F-sRRR4
RPRRNNsHLRDCCRGbRRRRRRRRR:RRRaQh )t ;-RR-GR bCFMMR0
RPRRNNsHLRDCCFGbMN_L#RCRR:RRRaQh )t ;-RR-GRCbCFMMF0RVCV#0R
RRNRPsLHNDVCRsRNORRRRRRRRRRR:)p qRRRR:j=R3Rj;RRRRR-R-RNwsOF0HMR
RRNRPsLHNDPCRN8DHVRbRRRRRRRR:PHND8b_V#00NCR;RRRRRR-R-RDeNHw8Ru0R#N
0CRRRRPHNsNCLDRbCGFRMRRRRRRRRR:hRz1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj
RRRR:RR=FR50sEC#>R=R''42R;RRRRRRRRRRRRRRR--e0COFxsHCC8RGMbFC
M0RCRLo
HMRRRRPHND8RVb:O=RD#N#V5bRN,soRCOEOC	_sssF2R;
RORRD#N#OCN#RO:RNR#CPHND8RVbHR#
RRRRRCIEM#RHGRR|b_F#xFCsRM|RCxo_CRsF|NRMMRR|JCkH0N_MM>R=
RRRRRRRR0sCkRsMj;3j
RRRRIRRERCMM_CoHRMV=R>
RRRRRsRRCs0kM R)qDp'FRI;RRRRRRRRRRRRR-RR-CRhoHN0PHCRMMVHH30$
RRRRIRRERCMb_F#HRMV=R>
RRRRRsRRCs0kM R)qEp'H;oERRRRRRRRRRRRR-RR-FRu#HH0PHCRMMVHH
0$RRRRRERICFMR0sEC#>R=
RRRRRRRRbCGFLM_NR#C:.=R*C*5GMbFC_M0I0H8E2-4R;-4
RRRRRRRRRHV0XF_jN45sCo5GMbFC_M0I0H8ER22=jR''ER0CRM
RRRRRRRRRo#HM=R:Rj43;R
RRRRRRDRC#RC
RRRRRRRRRo#HM=R:R3-4jR;
RRRRRCRRMH8RVR;
RRRRR-RR-HRwoCksR0FkRC0ERNVsOF0HMR
RRRRRRFRVsRRHHjMRRR0FVOsN0MHF_8IH04E-RFDFbR
RRRRRRRRRH0VRFj_X4s5No-R54RR-HR22=4R''ER0CRM
RRRRRRRRRVRRsRNO:V=RsRNO+.R53*jR*45-RH-R2
2;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8FRDFRb;RR--HR
RRRRRRVRHRDPNHb8VRb=RFM#_FNslDsRFRDPNHb8VRM=RCMo_FNslDsRFR0MFRM8CFNslDCHxRC0EMR
RRRRRRRRR-C-RGMbFCRM0/'=RjR',MlFsNVDRD0FNHRMobMFH0R
RRRRRRRRRCFGbMRRRRRRRRRRRRRRRRRRR:z=Rht1Qh5 7NRso5bCGFMMC0H_I8-0E4FR8IFM0R2j2;R
RRRRRRRRRCFGbMG5CbCFMMI0_HE80-R42:M=RFC0RGMbF5bCGFMMC0H_I8-0E4
2;RRRRRRRRRGRCbRRRRRRRRRRRRRRRRRRRR=R:R_0FHCM0oRCs5t1Qh5 7CFGbMR22+
4;RRRRRRRRRHR#oRMRRRRRRRRRRRRRRRRRR=R:Ro#HMRR*5j.3RR**C2GbR5*R4R3j+sRVN;O2
RRRRRRRR#CDC-RR-GRCbCFMM=0RR''j, RQ C RGM0C8RC8VNDF0oHMRHbFMR0
RRRRRRRRRbCGR=R:R-4RRbCGFLM_N;#C
RRRRRRRR#RRHRoM:#=RHRoM*.R53*jR*GRCb*2RRNVsOR;
RRRRRCRRMH8RVR;
RRRRRsRRCs0kMHR#o
M;RRRRCRM8OCN#RNOD#N#O#
C;RMRC8kRVMHO0F0MRFC_sN
D;
-RR-FRwsCResFHDoFROl0bNNDLHH
0$RkRVMHO0FsMRC0NDF0LH#NR5s:oRRq) ps2RCs0kMaR17p_zmBtQ_Be aRm)HR#
RPRRNNsHLRDCskC#D:0RRFVDNc0n;RRRRRRRR-RR-cRnR0LHRFVDNM0HoFRbH
M0RCRLo
HMRRRRskC#D:0R=FR0_FVDN50RNRso=N>Rs
o,RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>DRVFnN0cH'Eo
E,RRRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>VR-D0FNnDc'F;I2
RRRR0sCkRsM0#F_kRDP5#sCk2D0;R
RCRM8VOkM0MHFRNsCDL0FH;0#
R
RVOkM0MHFR0LH#s0FCRND5oNsR1:Raz7_pQmtB _eB)am2CRs0MksRq) p#RH
RRRRsPNHDNLCsRNoRnc:DRVFnN0cR;RRRRRRRRRRR--NRsoOPFMCCs08FR0RFVDNR0
RoLCHRM
RNRRsconRR:=0VF_D0FNRs5No>R=RoNs,R
RRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=V>RD0FNnEc'H,oE
RRRRRRRRRRRRRRRRRRRRRRRVOsN0MHF_8IH0=ER>VR-D0FNnDc'F;I2
RRRR0sCkRsM0sF_CRND5oNsn;c2
CRRMV8Rk0MOHRFML#H00CFsN
D;
-RR-kRbs#bFC):RCPlFCl#RC-0NDHFoORNDPkNDCV#RsRFlw#uR0MsHoR
RVOkM0MHFR_0Fj54R
RRRRoNsRRR:z h)1emp V7_D0FN;RRRRRRRRRRRRR--VNDF0oHMRHbFMH0RM0bk
RRRRqXvuRR:1_a7pQmtB=R:R''j2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0NR5sso'NCMo2R;
RoLCHRMR-V-Rk0MOHRFM0jF_4R
RRVRHRs5NoC'DMEo0R4<R2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRRRRR&"_amjR4:MDkDR08CCCO08s,RCs0kMoHMRphzpR"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRRsRRCs0kMqRhw
u;RRRRCRM8H
V;RRRRskC#D:0R=hRz)m 1p7e _FVDN50R1_a7pQmtB _eB)am5_0Fjz45ht1Qh5 70#F_DNP5s2o2,vRXq2u22R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFR_0Fj
4;
VRRk0MOHRFMQX#_
RRRRs5NoRR:z h)1emp V7_D0FN2R
RRCRs0MksRmAmph qR
H#RCRLo
HMRRRRskC0sQMR#R_X5_0F#5DPN2so2R;
R8CMRMVkOF0HM#RQ_
X;
VRRk0MOHRFM0XF_j54RNRso:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0NR5sso'NCMo2R;
RoLCHRM
RHRRVNR5sDo'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsw0Rpamq_ht  B)Q_tui'#HM0ONMCN_MlRC
RRRRR&RRRm"a_4Xj:kRMD8DRCO0C0,C8R0sCkHsMMhoRz"pp
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMhuqw;R
RRDRC#RC
RRRRR#sCkRD0:z=Rh1) m pe7D_VFRN05_0FX5j40#F_DNP5s2o22R;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0F0MRFj_X4
;
RkRVMHO0F0MRFj_X45ZRNRso:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0NR5sso'NCMo2R;
RoLCHRM
RHRRVNR5sDo'C0MoERR<402RE
CMRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRsFCbsw0Rpamq_ht  B)Q_tui'#HM0ONMCN_MlRC
RRRRR&RRRm"a_4XjZM:RkRDD8CC0O80C,CRs0MksHRMohpzp"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRRCRs0MksRwhquR;
RCRRD
#CRRRRRCRs#0kDRR:=z h)1emp V7_D0FNRF50_4XjZF50_P#D5oNs2;22
RRRRsRRCs0kMCRs#0kD;R
RRMRC8VRH;R
RCRM8VOkM0MHFR_0FXZj4;R

RMVkOF0HMFR0_jzX4NR5s:oRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNRs5NoN'sM2oC;R
RLHCoMR
RRVRHRs5NoC'DMEo0R4<R2ER0CRM
RRRRR#N#CRs0hWm_qQ)hhRt
RRRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRRRRR&"_amz4Xj:kRMD8DRCO0C0,C8R0sCkHsMMhoRz"pp
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR0sCkRsMhuqw;R
RRDRC#RC
RRRRR#sCkRD0:z=Rh1) m pe7D_VFRN05_0Fz4Xj5_0F#5DPN2so2
2;RRRRRCRs0MksR#sCk;D0
RRRR8CMR;HV
CRRMV8Rk0MOHRFM0zF_X;j4
R
R-a-RECC#RDNDFRI#0RECLCN#R0lNEkRVMHO0FRM#0kFR#0CRE8CRCkVNDP0RNCDk#R
R-F-RVER0CRHsbNNslCC0sR#3RkaE#ER0C8$RFkRVDQDR R  VNDF0oHMRHbFM
03RkRVMHO0F"MR+5"RDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sNMR858RDs,R2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR-5"RDs,RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0s#MRksL0NRO05RD,s
2;RMRC8kRVMHO0F"MR-
";
VRRk0MOHRFM"R*"5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
LRRCMoH
RRRR0sCkRsMl0kDH$bDR,5DR;s2
CRRMV8Rk0MOHRFM";*"
R
RVOkM0MHFR""/R,5DR:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RLHCoMR
RRCRs0MksRP8HHR8C5RD,s
2;RMRC8kRVMHO0F"MR/
";
VRRk0MOHRFM"lsC"DR5,RRs:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kMCRslMNH8RCs5RD,s
2;RMRC8kRVMHO0F"MRs"Cl;R

RMVkOF0HMlR"FR8"5RD,sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
LRRCMoH
RRRR0sCkRsMlkF8D5FRDs,R2R;
R8CMRMVkOF0HMlR"F;8"
R
R-F-RPDCsFCN88CRPsF#HMR#
RMVkOF0HM+R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR8N8R,5DRVs_D0FN2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"RDRR:)p q;RRs:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0,5DREs'H,oER'-sD2FI;R
RRCRs0MksR8N8R_5DVNDF0s,R2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR8N8R,5DRVs_D0FN2R;
R8CMRMVkOF0HM+R""
;
RkRVMHO0F"MR+5"RDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FN5RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMNR885VD_D0FN,2Rs;R
RCRM8VOkM0MHFR""+;R

RMVkOF0HM-R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRL#k0OsN0DR5,_RsVNDF0
2;RMRC8kRVMHO0F"MR-
";
VRRk0MOHRFM"R-"5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMkR#LN0sO50RDD_VF,N0R;s2
CRRMV8Rk0MOHRFM";-"
R
RVOkM0MHFR""-RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0s#MRksL0NRO05RD,sD_VF2N0;R
RCRM8VOkM0MHFR""-;R

RMVkOF0HM-R""DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0s#MRksL0NRO05VD_D0FN,2Rs;R
RCRM8VOkM0MHFR""-;R

RMVkOF0HM*R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRDlk0DHb$DR5,_RsVNDF0
2;RMRC8kRVMHO0F"MR*
";
VRRk0MOHRFM"R*"5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMkRlDb0HD5$RDD_VF,N0R;s2
CRRMV8Rk0MOHRFM";*"
R
RVOkM0MHFR""*RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0slMRkHD0bRD$5RD,sD_VF2N0;R
RCRM8VOkM0MHFR""*;R

RMVkOF0HM*R""DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0slMRkHD0bRD$5VD_D0FN,2Rs;R
RCRM8VOkM0MHFR""*;R

RMVkOF0HM/R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRP8HHR8C5RD,sD_VF2N0;R
RCRM8VOkM0MHFR""/;R

RMVkOF0HM/R""DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FN5RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsM8HHP85CRDD_VF,N0R;s2
CRRMV8Rk0MOHRFM";/"
R
RVOkM0MHFR""/RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0s8MRH8PHCDR5,_RsVNDF0
2;RMRC8kRVMHO0F"MR/
";
VRRk0MOHRFM"R/"5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0,5DREs'H,oER'-sD2FI;R
RRCRs0MksRP8HHR8C5VD_D0FN,2Rs;R
RCRM8VOkM0MHFR""/;R

RMVkOF0HMsR"CRl"5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpR0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0ssMRCHlNMs8CR,5DRVs_D0FN2R;
R8CMRMVkOF0HMsR"C;l"
R
RVOkM0MHFRC"sl5"RDRR:)p q;RRs:hRz)m 1p7e _FVDNR02skC0szMRh1) m pe7D_VFRN0HR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0,5DREs'H,oER'-sD2FI;R
RRCRs0MksRlsCN8HMC5sRDD_VF,N0R;s2
CRRMV8Rk0MOHRFM"lsC"
;
RkRVMHO0F"MRs"ClRR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0ssMRCHlNMs8CR,5DRVs_D0FN2R;
R8CMRMVkOF0HMsR"C;l"
R
RVOkM0MHFRC"sl5"RDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FN5RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMsNClHCM8sDR5_FVDNR0,s
2;RMRC8kRVMHO0F"MRs"Cl;R

RMVkOF0HMlR"FR8"5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpR0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0slMRFD8kFDR5,_RsVNDF0
2;RMRC8kRVMHO0F"MRl"F8;R

RMVkOF0HMlR"FR8"5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMFRl8FkDR_5DVNDF0s,R2R;
R8CMRMVkOF0HMlR"F;8"
R
RVOkM0MHFRF"l85"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR8lFkRDF5RD,sD_VF2N0;R
RCRM8VOkM0MHFRF"l8
";
VRRk0MOHRFM"8lF"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0slMRFD8kFDR5_FVDNR0,s
2;RMRC8kRVMHO0F"MRl"F8;R

RMVkOF0HM=R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMC5JRDs,R_FVDN;02
CRRMV8Rk0MOHRFM";="
R
RVOkM0MHFR="/"DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMM5CRDs,R_FVDN;02
CRRMV8Rk0MOHRFM""/=;R

RMVkOF0HM>R"=5"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2skC0sAMRm mpqHhR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRRoC5RD,sD_VF2N0;R
RCRM8VOkM0MHFR=">"
;
RkRVMHO0F"MR<R="5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpR0sCkRsMApmm RqhHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kMCRDR,5DRVs_D0FN2R;
R8CMRMVkOF0HM<R"=
";
VRRk0MOHRFM"R>"5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpR0sCkRsMApmm RqhHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kM0RoR,5DRVs_D0FN2R;
R8CMRMVkOF0HM>R""
;
RkRVMHO0F"MR<5"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2skC0sAMRm mpqHhR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRRD05RD,sD_VF2N0;R
RCRM8VOkM0MHFR""<;R

RMVkOF0HM=R""DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0sCMRJDR5_FVDNR0,s
2;RMRC8kRVMHO0F"MR=
";
VRRk0MOHRFM""/=RR5D: R)qRp;sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMCRMR_5DVNDF0s,R2R;
R8CMRMVkOF0HM/R"=
";
VRRk0MOHRFM"">=RR5D: R)qRp;sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMCRoR_5DVNDF0s,R2R;
R8CMRMVkOF0HM>R"=
";
VRRk0MOHRFM""<=RR5D: R)qRp;sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMCRDR_5DVNDF0s,R2R;
R8CMRMVkOF0HM<R"=
";
VRRk0MOHRFM"R>"5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm RqhHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0,5DREs'H,oER'-sD2FI;R
RRCRs0MksRRo05VD_D0FN,2Rs;R
RCRM8VOkM0MHFR"">;R

RMVkOF0HM<R""DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0sDMR0DR5_FVDNR0,s
2;RMRC8kRVMHO0F"MR<
";
VRRk0MOHRFM"R="5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  R)2skC0sAMRm mpqHhR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRRCJ5RD,sD_VF2N0;R
RCRM8VOkM0MHFR""=;R

RMVkOF0HM/R"=5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMM5CRDs,R_FVDN;02
CRRMV8Rk0MOHRFM""/=;R

RMVkOF0HM>R"=5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMo5CRDs,R_FVDN;02
CRRMV8Rk0MOHRFM"">=;R

RMVkOF0HM<R"=5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMD5CRDs,R_FVDN;02
CRRMV8Rk0MOHRFM""<=;R

RMVkOF0HM>R""DR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0soMR0DR5,_RsVNDF0
2;RMRC8kRVMHO0F"MR>
";
VRRk0MOHRFM"R<"5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  R)2skC0sAMRm mpqHhR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRRD05RD,sD_VF2N0;R
RCRM8VOkM0MHFR""<;R

RMVkOF0HM=R""DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMJRCR_5DVNDF0s,R2R;
R8CMRMVkOF0HM=R""
;
RkRVMHO0F"MR/R="5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpqHhR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FN5RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMM5CRDD_VF,N0R;s2
CRRMV8Rk0MOHRFM""/=;R

RMVkOF0HM>R"=5"RDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMmRAmqp h#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VF5N0Ds,R'oEHE-,RsF'DI
2;RRRRskC0soMRCDR5_FVDNR0,s
2;RMRC8kRVMHO0F"MR>;="
R
RVOkM0MHFR="<"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksRmAmph qR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDND05,'RsEEHo,sR-'IDF2R;
RsRRCs0kMCRDR_5DVNDF0s,R2R;
R8CMRMVkOF0HM<R"=
";
VRRk0MOHRFM"R>"5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0sAMRm mpqHhR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FN5RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMo50RDD_VF,N0R;s2
CRRMV8Rk0MOHRFM";>"
R
RVOkM0MHFR""<RR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsMApmm RqhHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0,5DREs'H,oER'-sD2FI;R
RRCRs0MksRRD05VD_D0FN,2Rs;R
RCRM8VOkM0MHFR""<;R

RR--?F=RPDCsF#N8
VRRk0MOHRFM""?=RR5D:hRz)m 1p7e _FVDNR0;sRR:)p q2CRs0MksR71a_mzptRQBHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kMRRD?s=R_FVDN
0;RMRC8kRVMHO0F"MR?;="
R
RVOkM0MHFR/"?=5"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMD/R?=_RsVNDF0R;
R8CMRMVkOF0HM?R"/;="
R
RVOkM0MHFR>"?"DR5Rz:Rh1) m pe7D_VF;N0R:sRRq) ps2RCs0kMaR17p_zmBtQR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0sDMRRR?>sD_VF;N0
CRRMV8Rk0MOHRFM""?>;R

RMVkOF0HM?R">R="5:DRR)zh p1me_ 7VNDF0s;RR):R 2qpR0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR?DR>s=R_FVDN
0;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<5"RDRR:z h)1emp V7_D0FN;RRs: R)qRp2skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMD<R?RVs_D0FN;R
RCRM8VOkM0MHFR<"?"
;
RkRVMHO0F"MR?"<=RR5D:hRz)m 1p7e _FVDNR0;sRR:)p q2CRs0MksR71a_mzptRQBHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kMRRD?R<=sD_VF;N0
CRRMV8Rk0MOHRFM"=?<"
;
R-R-RNsCDMRN8DRVF
N0RkRVMHO0F"MR?R="5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FNR,5DREs'H,oER'-sD2FI;R
RRCRs0MksRVD_D0FNRR?=sR;
R8CMRMVkOF0HM?R"=
";
VRRk0MOHRFM"=?/"DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0s2RCs0kMaR17p_zmBtQR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDN50RDs,R'oEHE-,RsF'DI
2;RRRRskC0sDMR_FVDN?0R/s=R;R
RCRM8VOkM0MHFR/"?=
";
VRRk0MOHRFM""?>RR5D: R)qRp;sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzptRQBHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0DR5,'RsEEHo,sR-'IDF2R;
RsRRCs0kM_RDVNDF0>R?R
s;RMRC8kRVMHO0F"MR?;>"
R
RVOkM0MHFR>"?=5"RDRR:)p q;RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VFRN05RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMDD_VFRN0?R>=sR;
R8CMRMVkOF0HM?R">;="
R
RVOkM0MHFR<"?"DR5R):R ;qpR:sRR)zh p1me_ 7VNDF0s2RCs0kMaR17p_zmBtQR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDN50RDs,R'oEHE-,RsF'DI
2;RRRRskC0sDMR_FVDN?0R<;Rs
CRRMV8Rk0MOHRFM""?<;R

RMVkOF0HM?R"<R="5:DRRq) ps;RRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FNR,5DREs'H,oER'-sD2FI;R
RRCRs0MksRVD_D0FNR=?<R
s;RMRC8kRVMHO0F"MR?"<=;R

RR--?F=RPDCsF#N8
VRRk0MOHRFM""?=RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR?DR=_RsVNDF0R;
R8CMRMVkOF0HM?R"=
";
VRRk0MOHRFM"=?/"DR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2CRs0MksR71a_mzptRQBHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kMRRD?R/=sD_VF;N0
CRRMV8Rk0MOHRFM"=?/"
;
RkRVMHO0F"MR?R>"5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  R)2skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMD>R?RVs_D0FN;R
RCRM8VOkM0MHFR>"?"
;
RkRVMHO0F"MR?">=RR5D:hRz)m 1p7e _FVDNR0;sRR:Q hat2 )R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksR?DR>s=R_FVDN
0;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<5"RDRR:z h)1emp V7_D0FN;RRs:hRQa  t)s2RCs0kMaR17p_zmBtQR
H#RRRRPHNsNCLDRVs_D0FNRz:Rh1) m pe7D_VFRN05sD'NCMo2R;
RoLCHRM
RsRR_FVDN:0R=FR0_FVDN50RsD,R'oEHE-,RDF'DI
2;RRRRskC0sDMRRR?<sD_VF;N0
CRRMV8Rk0MOHRFM""?<;R

RMVkOF0HM?R"<R="5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  R)2skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMD<R?=_RsVNDF0R;
R8CMRMVkOF0HM?R"<;="
R
R-H-RMo0CCNsRMV8RD0FN
VRRk0MOHRFM""?=RR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FNR,5DREs'H,oER'-sD2FI;R
RRCRs0MksRVD_D0FNRR?=sR;
R8CMRMVkOF0HM?R"=
";
VRRk0MOHRFM"=?/"DR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2CRs0MksR71a_mzptRQBHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0DR5,'RsEEHo,sR-'IDF2R;
RsRRCs0kM_RDVNDF0/R?=;Rs
CRRMV8Rk0MOHRFM"=?/"
;
RkRVMHO0F"MR?R>"5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VFRN05RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMDD_VFRN0?s>R;R
RCRM8VOkM0MHFR>"?"
;
RkRVMHO0F"MR?">=RR5D:hRQa  t)s;RRz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RRNRPsLHNDDCR_FVDN:0RR)zh p1me_ 7VNDF0sR5'MsNo;C2
LRRCMoH
RRRRVD_D0FNRR:=0VF_D0FNR,5DREs'H,oER'-sD2FI;R
RRCRs0MksRVD_D0FNR=?>R
s;RMRC8kRVMHO0F"MR?">=;R

RMVkOF0HM?R"<5"RDRR:Q hat; )R:sRR)zh p1me_ 7VNDF0s2RCs0kMaR17p_zmBtQR
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDN50RDs,R'oEHE-,RsF'DI
2;RRRRskC0sDMR_FVDN?0R<;Rs
CRRMV8Rk0MOHRFM""?<;R

RMVkOF0HM?R"<R="5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VFRN05RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMDD_VFRN0?R<=sR;
R8CMRMVkOF0HM?R"<;="
R
R-l-RHlMHkNlRMl8RNlGHkFlRPDCsF#N8
VRRk0MOHRFMlHHMlRkl5:DRR)zh p1me_ 7VNDF0s;RR):R 2qp
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCR_FVDN:0RR)zh p1me_ 7VNDF0DR5'MsNo;C2
LRRCMoH
RRRRVs_D0FNRR:=0VF_D0FNR,5sRED'H,oER'-DD2FI;R
RRCRs0MksRMlHHllkR,5DRVs_D0FN2R;
R8CMRMVkOF0HMHRlMkHll
;
RkRVMHO0FlMRNlGHk5lRDRR:z h)1emp V7_D0FN;RRs: R)q
p2RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMlHNGlRkl5RD,sD_VF2N0;R
RCRM8VOkM0MHFRGlNHllk;R

RMVkOF0HMHRlMkHllDR5R):R ;qpR:sRR)zh p1me_ 7VNDF0R2
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDRVD_D0FNRz:Rh1) m pe7D_VFRN05ss'NCMo2R;
RoLCHRM
RDRR_FVDN:0R=FR0_FVDN50RDs,R'oEHE-,RsF'DI
2;RRRRskC0slMRHlMHk5lRDD_VF,N0R;s2
CRRMV8Rk0MOHRFMlHHMl;kl
R
RVOkM0MHFRGlNHllkRR5D: R)qRp;sRR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0DR5,'RsEEHo,sR-'IDF2R;
RsRRCs0kMNRlGkHllDR5_FVDNR0,s
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5:DRR)zh p1me_ 7VNDF0s;RRQ:Rhta  
)2RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLC_RsVNDF0RR:z h)1emp V7_D0FNR'5DsoNMC
2;RCRLo
HMRRRRsD_VFRN0:0=RFD_VFRN05Rs,DH'EoRE,-DD'F;I2
RRRR0sCkRsMlHHMlRkl5RD,sD_VF2N0;R
RCRM8VOkM0MHFRMlHHllk;R

RMVkOF0HMNRlGkHllDR5Rz:Rh1) m pe7D_VF;N0R:sRRaQh )t 2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCsD_VFRN0:hRz)m 1p7e _FVDN50RDN'sM2oC;R
RLHCoMR
RR_RsVNDF0=R:R_0FVNDF0sR5,'RDEEHo,DR-'IDF2R;
RsRRCs0kMNRlGkHllDR5,_RsVNDF0
2;RMRC8kRVMHO0FlMRNlGHk
l;
VRRk0MOHRFMlHHMlRkl5:DRRaQh )t ;RRs:hRz)m 1p7e _FVDN
02RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLC_RDVNDF0RR:z h)1emp V7_D0FNR'5ssoNMC
2;RCRLo
HMRRRRDD_VFRN0:0=RFD_VFRN05RD,sH'EoRE,-Ds'F;I2
RRRR0sCkRsMlHHMlRkl5VD_D0FN,2Rs;R
RCRM8VOkM0MHFRMlHHllk;R

RMVkOF0HMNRlGkHllDR5RQ:Rhta  R);sRR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCDD_VFRN0:hRz)m 1p7e _FVDN50RsN'sM2oC;R
RLHCoMR
RR_RDVNDF0=R:R_0FVNDF0DR5,'RsEEHo,sR-'IDF2R;
RsRRCs0kMNRlGkHllDR5_FVDNR0,s
2;RMRC8kRVMHO0FlMRNlGHk
l;
-RR-------------------------------------------------------------------------
--R-R-RoDFHDONRMVkOF0HMR#
R----------------------------------------------------------------------------R
RVOkM0MHFRF"M05"RpRR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC R)1azpR1:Raz7_pQmtB _eB)am5Dp'C0MoER-48MFI0jFR2R;R-V-RFCsORI8FM
0FRCRLo
HMRRRR)z 1p:aR=FRM0FR0_D#kP25p;R
RRCRs0MksR_0FVNDF0)R5 p1zap,R'oEHE-,RpF'DI
2;RMRC8kRVMHO0F"MRM"F0;R

RMVkOF0HMNR"MR8"5Rp,)RR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC R)1azpR1:Raz7_pQmtB _eB)am5Dp'C0MoER-48MFI0jFR2R;R-V-RFCsORI8FM
0FRLRRCMoH
RRRRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pR8NMR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"M"N8:""RM)NoCCRsssFR)p'q htRR/=)q')h"t 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR1) zRpa:5=RFC0Es=#R>XR''
2;RRRRCRM8H
V;RRRRskC0s0MRFD_VFRN051) z,paREp'H,oER'-pD2FI;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM""FsR,5pR:)RR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHND)CR p1zaRR:1_a7ztpmQeB_ mBa)'5pDoCM04E-RI8FMR0FjR2;RR--VOFsCFR8IFM0
LRRCMoH
RRRRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRRFs0#F_k5DP)
2;RRRRCCD#
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRR&"R"""Fs"):RNCMoRsCsFpsR'h)qt/ R='R))tqh R"
RRRRR#RRCsPCHR0$IMNsH;Mo
RRRR)RR p1za=R:R05FE#CsRR=>'2X';R
RRMRC8VRH;R
RRCRs0MksR_0FVNDF0)R5 p1zap,R'oEHE-,RpF'DI
2;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRN"MMR8"5Rp,)RR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC R)1azpR1:Raz7_pQmtB _eB)am5Dp'C0MoER-48MFI0jFR2R;R-V-RFCsORI8FM
0FRCRLo
HMRRRRRRHV5Ep'HRoE='R)EEHoR8NMRDp'F=IRRD)'FRI20MEC
RRRR)RR p1za=R:R_0F#PkD5Rp2M8NMR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"N"MM"8":NR)MRoCCFsss'Rp)tqh =R/R))'q ht"R
RRRRRRCR#PHCs0I$RNHsMM
o;RRRRR R)1azpRR:=5EF0CRs#='>RX;'2
RRRR8CMR;HV
RRRR0sCkRsM0VF_D0FNR 5)1azp,'RpEEHo,pR-'IDF2R;
R8CMRMVkOF0HMMR"N"M8;R

RMVkOF0HMMR"FRs"5Rp,)RR:z h)1emp V7_D0FN2CRs0MksR)zh p1me_ 7VNDF0#RH
RRRRsPNHDNLC R)1azpR1:Raz7_pQmtB _eB)am5Dp'C0MoER-48MFI0jFR2R;R-V-RFCsORI8FM
0FRCRLo
HMRRRRRRHV5Ep'HRoE='R)EEHoR8NMRDp'F=IRRD)'FRI20MEC
RRRR)RR p1za=R:R_0F#PkD5Rp2MRFs0#F_k5DP)
2;RRRRCCD#
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""sMF"R":)oNMCsRCsRFspq')hRt /)=R'h)qt
 "RRRRRRRR#CCPs$H0RsINMoHM;R
RRRRR)z 1p:aR=FR50sEC#>R=R''X2R;
RCRRMH8RVR;
RsRRCs0kMFR0_FVDN50R)z 1pRa,pH'EoRE,-Dp'F;I2
CRRMV8Rk0MOHRFM"sMF"
;
RkRVMHO0F"MRG"FsR,5pR:)RR)zh p1me_ 7VNDF0s2RCs0kMhRz)m 1p7e _FVDNH0R#R
RRNRPsLHND)CR p1zaRR:1_a7ztpmQeB_ mBa)'5pDoCM04E-RI8FMR0FjR2;RR--VOFsCFR8IFM0
LRRCMoH
RRRRVRHR'5pEEHoR)=R'oEHEMRN8'RpDRFI='R)D2FIRC0EMR
RRRRR)z 1p:aR=FR0_D#kP25pRsGFR_0F#PkD5;)2
RRRR#CDCR
RRRRRNC##sh0Rmq_W)hhQtR
RRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNl
RRRRRRRR"&R"F"Gs:""RM)NoCCRsssFR)p'q htRR/=)q')h"t 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR1) zRpa:5=RFC0Es=#R>XR''
2;RRRRCRM8H
V;RRRRskC0s0MRFD_VFRN051) z,paREp'H,oER'-pD2FI;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"Rp),RRz:Rh1) m pe7D_VF2N0R0sCkRsMz h)1emp V7_D0FNR
H#RRRRPHNsNCLDR1) zRpa:aR17p_zmBtQ_Be a5m)pC'DMEo0-84RF0IMF2Rj;-RR-FRVsROC8MFI0RF
RoLCHRM
RRRRH5VRpH'Eo=ERRE)'HRoENRM8pF'DIRR=)F'DI02RE
CMRRRRR R)1azpRR:=0#F_k5DPpG2RMRFs0#F_k5DP)
2;RRRRCCD#
RRRRNRR#s#C0mRh_)WqhtQh
RRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRR&"R""FGMs:""RM)NoCCRsssFR)p'q htRR/=)q')h"t 
RRRRRRRRP#CC0sH$NRIsMMHoR;
RRRRR1) zRpa:5=RFC0Es=#R>XR''
2;RRRRCRM8H
V;RRRRskC0s0MRFD_VFRN051) z,paREp'H,oER'-pD2FI;R
RCRM8VOkM0MHFRM"GF;s"
R
R-e-RCFO0sMRN80R#8D_kFOoHRMVkOF0HMR#,#CNlRRN#VOkM0MHF#MRHRlMkCOsH_8#0
VRRk0MOHRFM"8NM"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7D_VF2N0
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5)soNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50RpMRN8FR0_D#kP25)2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM"8NM"pR5Rz:Rh1) m pe7D_VF;N0R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5psoNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50R0#F_k5DPpN2RM)8R2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRM"N8
";
VRRk0MOHRFM""FsRR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _FVDN
02RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7D_VFRN05s)'NCMo2R;
RoLCHRM
RsRRCD#k0=R:R)zh p1me_ 7VNDF0pR5RRFs0#F_k5DP);22
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRF;s"
R
RVOkM0MHFRs"F"pR5Rz:Rh1) m pe7D_VF;N0R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5psoNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50R0#F_k5DPpF2Rs2R);R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM""Fs;R

RMVkOF0HMMR"N"M8RR5p:aR17p_zmBtQ;RR):hRz)m 1p7e _FVDN
02RRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRsPNHDNLCCRs#0kDRz:Rh1) m pe7D_VFRN05s)'NCMo2R;
RoLCHRM
RsRRCD#k0=R:R)zh p1me_ 7VNDF0pR5RMMN8FR0_D#kP25)2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRN"MM;8"
R
RVOkM0MHFRN"MMR8"5:pRR)zh p1me_ 7VNDF0);RR1:Raz7_pQmtBR2
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _FVDN50RpN'sM2oC;R
RLHCoMR
RRCRs#0kDRR:=z h)1emp V7_D0FNRF50_D#kP25pRMMN82R);R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFM"MMN8
";
VRRk0MOHRFM"sMF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7D_VF2N0
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5)soNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50RpFRMsFR0_D#kP25)2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Ms
";
VRRk0MOHRFM"sMF"pR5Rz:Rh1) m pe7D_VF;N0R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5psoNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50R0#F_k5DPpM2RF)sR2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Ms
";
VRRk0MOHRFM"sGF"pR5R1:Raz7_pQmtB);RRz:Rh1) m pe7D_VF2N0
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5)soNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50RpFRGsFR0_D#kP25)2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"sGF"pR5Rz:Rh1) m pe7D_VF;N0R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5psoNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50R0#F_k5DPpG2RF)sR2R;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRF"Gs
";
VRRk0MOHRFM"FGMs5"RpRR:1_a7ztpmQRB;)RR:z h)1emp V7_D0FN2R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0)R5'MsNo;C2
LRRCMoH
RRRR#sCkRD0:z=Rh1) m pe7D_VFRN05GpRMRFs0#F_k5DP);22
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0F"MRGsMF"
;
RkRVMHO0F"MRGsMF"pR5Rz:Rh1) m pe7D_VF;N0R:)RR71a_mzpt2QB
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNR'5psoNMC
2;RCRLo
HMRRRRskC#D:0R=hRz)m 1p7e _FVDN50R0#F_k5DPpG2RMRFs)
2;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMGR"M"Fs;R

RR--)kC8OF0HMbRFC0sNF,s#Rl#NC#RNRlMkCOsH_8#0RMVkOF0HM
#
RkRVMHO0F"MRN"M8RR5D:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMNRM80#F_k5DPD
2;RMRC8kRVMHO0F"MRN"M8;R

RMVkOF0HMMR"N"M8RR5D:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMM8NMR_0F#PkD5;D2
CRRMV8Rk0MOHRFM"MMN8
";
VRRk0MOHRFM""FsRR5D:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMF0sRFk_#DDP52R;
R8CMRMVkOF0HMFR"s
";
VRRk0MOHRFM"sMF"DR5Rz:Rh1) m pe7D_VF2N0R0sCkRsM1_a7ztpmQHBR#R
RLHCoMR
RRCRs0MksRsMFR_0F#PkD5;D2
CRRMV8Rk0MOHRFM"sMF"
;
RkRVMHO0F"MRG"FsRR5D:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMGRFs0#F_k5DPD
2;RMRC8kRVMHO0F"MRG"Fs;R

RMVkOF0HMGR"M"FsRR5D:hRz)m 1p7e _FVDNR02skC0s1MRaz7_pQmtB#RH
LRRCMoH
RRRR0sCkRsMGsMFR_0F#PkD5;D2
CRRMV8Rk0MOHRFM"FGMs
";
-RR----------------------------------------------------------------------------
-RR-CR)OlFlCCM88kRwMHO0FRM#VlsFRC0ER Q  6R(cbRqb8CMHRG
R----------------------------------------------------------------------------R-
RR--skC0sRM#GHRI00ERE#CRHRoMF$VR3R
RVOkM0MHFRbBF$o#HM
R5RRRRG$,RRz:Rh1) m pe7D_VF2N0RRRRRRRRRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRskC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kM5R$$H'EoRE2&RRG5EG'H-oE4FR8IFM0RDG'F;I2
CRRMV8Rk0MOHRFMB$Fb#MHo;R

RR--)kC0sRM#$RR*.M**RsVFR0HMCNosDNRPD#kCRRFVhHRI0kEF0FROl0bkHRMo.M**
VRRk0MOHRFM1DONL
R5RRRR$RRRRRRRRRRRRRRRRRRRRz:Rh1) m pe7D_VF;N0RRRRR-R-RFVDNM0HoFRbHRM0HkMb0R
RRRRhRRRRRRRRRRRRRRRRR:RRRaQh )t ;RRRR-R-RbCGFMMC0FR0R8N8RRRR
RRRRMOF#M0N0FRsk_M8#D0$CRR:sMFk8$_0b:CR=DRVF_N0sMFk80_#$;DCR-R-RksFMM8HobRF0MHF
RRRRMOF#M0N0EROC_O	CFsssRR:Apmm RqhR:RR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRRRR:V=RD0FN_M8CFNslDCHx2-RR-#RzC RQ C RGM0C8RC8wRu
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RH-lM$C5'IDF,'R$D2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=$H'EoRE;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRsPNHDNLCsRNos,RCD#k0RRRRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0;E2R-R-R0HMCNsMDsRNoCklMR0
RPRRNNsHLRDCCFGbMRRRRRRRR:RRRt1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2R-R-ROeC0HFsxRC8C
GbRRRRPHNsNCLDRbCGRRRRRRRRRRRR:QR1t7h RG5CbCFMMI0_HE80RI8FMR0Fj
2;RRRRPHNsNCLDRskVNRO0RRRRRRRR:hRz1hQt 57RVOsN0MHF_8IH08ERF0IMF2Rj;R
RRFROMN#0MC0RGMbF_#LNCRRRRRR:1hQt 57RCFGbM0CM_8IH04E-RI8FMR0FjR2
RRRRRR:=o_CMCFGbMN_L#CC5GMbFC_M0I0H8ER2;RRRRRRRRRR--CFGbM0CMRVFV#
C0RRRRPHNsNCLDR0Vb$RbC:NRPD_H8V0b#N;0C
LRRCMoH
RRRRR--a#EHRMONRRLC8CFMRRL$#bHlDN$R8M8HoRRh00FRECCRGMbFC3M0
RRRRoNsRRRR:0=RF4_jR,5$R''X2R;
RVRRbb0$C=R:RNOD#b#V5oNs,EROC_O	CFsss
2;RRRRO#DN##ONCRR:OCN#R0Vb$RbCHR#
RRRRRCIEM#RHG>R=
RRRRRRRR#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRRERICMMRN|MRRHJkCM0_N=MR>R
RRRRRR-R-R0)CkRsMJCkH0qRhhQ,R (  64c-g-U6(,344R
RRRRRRCRs#0kDRR:=JMMNV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRCIEM0RFE#CsR
=>RRRRRRRRLNsC	k_MlsLCRR5
RRRRRRRRRoNsRRRRRRRRRR=>N,so
RRRRRRRRVRRbb0$RRRRR=RR>bRV0C$b,R
RRRRRRRRR8FCMsDlNHRxC=8>RCsMFlHNDx
C,RRRRRRRRRsRVNRO0RRRRR>R=RskVN,O0
RRRRRRRRCRRGMbFRRRRR=RR>GRCb2FM;R
RRRRRRGRCb=R:R#sCHRxC5bCGFRM,C'GbDoCM0RE2+;Rh
RRRRRRRR#sCkRD0:M=RFNslDCHxRR5
RRRRRRRRRNVsOR0RRRRRRRRR=k>RVOsN0R,
RRRRRRRRRbCGFRMRRRRRRRRR=C>RG
b,RRRRRRRRRHR#oRMRRRRRRRRRRR=>0GF_j54RNRso5oNs'oEHE,22
RRRRRRRRVRRs0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRCRRGMbFC_M0I0H8E>R=RbCGFMMC0H_I8,0E
RRRRRRRRsRRF8kM_$#0DRCRR>R=RksFM#8_0C$D,R
RRRRRRRRR8FCMsDlNHRxCR=RR>CR8MlFsNxDHCR,
RRRRRRRRRkMoNRs8RRRRRRRR=j>R2R;
RCRRMO8RNR#CO#DN##ONCR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRN1OD
L;
-RR-CR)0Mks#RR$**R.*VMRFHsRMo0CsRNDPkNDCF#RVRRhIEH0FRk0ObFlkM0Ho*R.*RM
RMVkOF0HMOR1NRDL5R
RRRR$RRRRRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRR--VNDF0oHMRHbFMH0RM0bk
RRRRRhRRRRRRRRRRRRRRRRRRRR:z h)1emp 17_Q th7R;R-C-RGMbFCRM00NFR8R8RRRR
RORRF0M#NRM0sMFk80_#$RDC:FRsk_M80C$bRR:=VNDF0F_sk_M8#D0$CR;R-s-RF8kMHRMoFHb0FRM
RORRF0M#NRM0OOEC	s_CsRFs:mRAmqp hRRRRR:=VNDF0E_OC_O	CFsssR;R-O-RE	CORsVFRsCsF
s#RRRRO#FM00NMRM8CFNslDCHxRA:Rm mpqRhRR=R:RFVDN80_CsMFlHNDxRC2RR--zR#CQ   R0CGCCM88uRw
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDMCR_0HMRQ:Rhta  
);RCRLo
HMRRRRMM_H0=R:R_0FHCM0o5Csh
2;RRRRskC0s1MROLNDRR5$RRRRRRRRR>R=R
$,RRRRRRRRRRRRRRRRRRRhRRRRRRRRR>R=RHM_M
0,RRRRRRRRRRRRRRRRRFRsk_M8#D0$C>R=RksFM#8_0C$D,R
RRRRRRRRRRRRRRRRROOEC	s_CsRFs=O>RE	CO_sCsF
s,RRRRRRRRRRRRRRRRRCR8MlFsNxDHC>R=RM8CFNslDCHx2R;
R8CMRMVkOF0HMOR1N;DL
R
R-s-RCs0kM0#REkCRMNLH#RC8CFGbM0CMRRFVGR
RVOkM0MHFRopFL
R5RRRRGRR:z h)1emp V7_D0FN2RRRRRRRRRRRRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRskC0sQMRhta  R)
R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RH-lM5CRGF'DIG,R'IDF2R;R-D-RC0MoEVRFRRwuFbk0kV0Rs0NOH
FMRRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:REG'H;oER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHNDsCRCD#k0RRRRRRRRRR:Q hat; )R-R-R#sCk
D0RRRRPHNsNCLDRoNsRRRRRRRRRRRR:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8ER2;RR--HCM0sDMNRoNskMlC0R
RRNRPsLHNDCCRGMbFRRRRRRRRRRR:1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj;R
RRNRPsLHNDVCRs0NORRRRRRRRRRR:zQh1t7h Rs5VNHO0FIM_HE80RI8FMR0Fj
2;RRRRO#FM00NMRbCGFLM_NR#CRRRR:hRQa  t)=R:R*.*5bCGFMMC0H_I8-0E4-2R4R;R-C-RGMbFC
M0RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-F-RVCV#04R+
RRRRsPNHDNLCbRV0C$bRRRRRRRRRP:RN8DH_#Vb0CN0;R
RLHCoMR
RR-R-R#Kk0CRs0MksRC0ERbCGFMMC0R3
RNRRsRoRR=R:R_0Fj54RG',RX;'2
RRRR0Vb$RbC:O=RD#N#VNb5s;o2
RRRRNOD#N#O#:CRR#ONCbRV0C$bR
H#RRRRRERICHMR#|GRRMMNRJ|Rk0HC_MMNR
=>RRRRRRRR-)-RCs0kMkRJHRC0h,qhR Q  c(6-U4g63-(4
,4RRRRRRRRskC#D:0R=;Rj
RRRRIRRERCMb_F#8FCMsDlNRM|RC8o_CsMFlRND=R>
RRRRRVRRs0NORs5VNHO0FIM_HE802=R:R''j;R
RRRRRRsRVNRO05NVsOF0HMH_I8-0E4FR8IFM0RRj2:R=
RRRRRRRRR1zhQ th70R5FD_#Ps5No45-RI8FMR0F-NVsOF0HMH_I820E2
2;RRRRRRRRskC#D:0R=HRVMD8_ClV0FR#05NVsOR0,'24'RRRRR-R-RMwH8ER0CHRVsR#0"
4"RRRRRRRRRRRRRRRRRRR-VOsN0MHF_8IH0RE;RRRR-#-RksL0NRO00RECDoCM0IERCNRIMR0
RRRRRsRRCD#k0=R:RG-Cb_FMLCN#R4+RRs+RCD#k0R;
RRRRRCIEM0RFE#CsR
=>RRRRRRRRCFGbMRRRRRRRRRRRRRRRRRRR:1=RQ th7s5NoCR5GMbFC_M0I0H8ERR-4FR8IFM0R2j2;R
RRRRRRGRCb5FMCFGbM0CM_8IH04E-2=R:R0MFRbCGFCM5GMbFC_M0I0H8E2-4;R
RRRRRRGRCbRFMRRRRRRRRRRRRRRRRR=R:RbCGF+MRR
4;RRRRRRRRskC#DR0RRRRRRRRRRRRRRRRR:0=RFM_H0CCosCR5GMbF2R;
RCRRMO8RNR#CO#DN##ONCR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRopFL
;
R-R-R0sCk#sMRC0ERLkMHCN#8GRCbCFMMF0RV
RGRkRVMHO0FpMRFRoL5R
RRRRG:hRz)m 1p7e _FVDNR02RRRRRRRRRRRRR-R-RFVDNM0HoFRbHRM0HkMb0R
RRCRs0MksR)zh p1me_ 71hQt R7
R
H#RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:REG'H;oER-R-RMDCoR0EFwVRukRF00bkRbCGFMMC0R
RRNRPsLHNDsCRCD#k0RRRRRRRRRR:1hQt 57RCFGbM0CM_8IH0-ERR84RF0IMF2Rj;-RR-CRs#0kD
LRRCMoH
RRRRR--K0k#R0sCkRsM0RECCFGbM0CM3R
RRCRs#0kDRR:=0#F_HCoM8pR5FRoL5,G2RbCGFMMC0H_I820E;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMpLFo;R

RR--skC0sRM#0RECM0CGRbsCsCC#ML0NDMCRCEHoLRFsFGVRRRHM0REC8CHsOF0HMFR0I8NsRR$
RMVkOF0HMCRhGV0N0RCs5R
RR,RGRR$RRRRRRRRRRRRRR:RRR)zh p1me_ 7VNDF0R;RRRRR-V-RD0FNHRMobMFH0MRHb
k0RRRRO#FM00NMRCOEOC	_sssFRA:Rm mpq:hR=DRVF_N0OOEC	s_Cs;FsR-R-RCOEOV	RFCsRsssF#R
RRFROMN#0M80RCsMFlHNDx:CRRmAmph qRR:=VNDF0C_8MlFsNxDHCR2
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RH-lMGC5'IDF,'RGD2FI;-RR-CRDMEo0RRFVwFuRkk0b0sRVNHO0FRM
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=GH'EoRE;RR--DoCM0FERVuRwR0FkbRk0CFGbM0CM
RRRRMVkOF0HM=R""
R5RRRRR,RDR:sRR)zh p1me_ 7VNDF0R2RRRRRRRRR-H-RM0bk#R
RRRRRskC0sAMRm mpqHhR#R
RRCRLoRHMRR--VOkM0MHFR""=
RRRRsRRCs0kMJRCRR5DRRRRRRRRR>R=R
D,RRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=>sR,
RRRRRRRRRRRRRRRROOEC	s_CsRFs=V>RNCD#2R;
RCRRMV8Rk0MOHRFM";="
RRRRMVkOF0HM>R""
R5RRRRR,RDR:sRR)zh p1me_ 7VNDF0R2RRRRRRRRR-H-RM0bk#R
RRRRRskC0sAMRm mpqHhR#R
RRCRLoRHMRR--VOkM0MHFR"">
RRRRsRRCs0kM0RoRR5DRRRRRRRRR>R=R
D,RRRRRRRRRRRRRRRRRRsRRRRRRRRRRR=>sR,
RRRRRRRRRRRRRRRROOEC	s_CsRFs=V>RNCD#2R;
RCRRMV8Rk0MOHRFM";>"
RRRRsPNHDNLCsRVNRO0RRRRRRRRRRRRRz:Rht1QhR 75NVsOF0HMH_I8-0E4FR8IFM0R;j2
RRRRsPNHDNLCGRCbRFMRRRRRRRRRRRRRz:Rht1QhR 75bCGFMMC0H_I8-0E4FR8IFM0R;j2
RRRRsPNHDNLCHR#oRMRRRRRRRRRRRRRR1:Raz7_pQmtBR;
RPRRNNsHLRDCskC#DR0RRRRRRRRRR:RRR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RPRRNNsHLRDCPHND8GVb,NRPDVH8b:$RRDPNHV8_bN#00RC;RR--eHND8uRwRN#00RC
RoLCHRMR-V-RbC_hGV0N0
CsRRRR-Q-RVRRY>,RXR8N8RCFMRR0F0RECVOsN0MHF,0RFEICsHR#C#0kLs0NO3R
RRNRPDVH8b:GR=DRONV##bGR5,EROC_O	CFsss
2;RRRRPHND8$VbRR:=O#DN#RVb5R$,OOEC	s_Cs2Fs;R
RRVRHRDPNHb8VGRR=HR#GFPsRN8DHVRb$=#RHGER0CRM
RRRRR#sCkRD0:5=RFC0Es=#R>XR''
2;RRRRRCRs0MksR#sCk;D0
RRRR#CDH5VRPHND8GVbRM=RNFMRsNRPDVH8b=$RRMMN2ER0CRM
RRRRR0sCkRsMMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRCHD#VPR5N8DHVRbG=kRJH_C0MRNMFPsRN8DHVRb$=kRJH_C0M2NMRC0EMR
RRRRRskC0sJMRMVNMbVR5s0NOH_FMI0H8E>R=RNVsOF0HMH_I8,0E
RRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRR#CDHGVRR$=RRC0EMRRRRRRRRRRRRRRRRRRRRR--)kC0sXMR
RRRRsRRCs0kM;RG
RRRR#CDCR
RRRRRVOsN0=R:R1zhQ th70R5FD_#PGR5R45-RI8FMR0F-NVsOF0HMH_I820E2R2;RR--wOsN0MHF
RRRRCRRGMbFRR:=zQh1t7h RR5G5bCGFMMC0H_I8R0E-RR48MFI0jFR2R2;RRRR-C-RGMbFC
M0RRRRRHR#oRMR:G=R5bCGFMMC0H_I820E;RRRRRRR-#-RHRoML
H0RRRRRVRHRR5$>2RGRC0EMR
RRRRRR-R-ROQMs#CNCER0CkRMlsLCRPoHCRM
RRRRRHRRVNRPDVH8b=GRRoMC_VHMRC0EMR
RRRRRRRRR-s-RCs0kMFRl#M0RC0oNHRPCMLklCRs
RRRRRRRRRbCGFRMRR:RR=FR50sEC#>R=R''42R;
RRRRRRRRRbCGF5MRj:2R=jR''R;
RRRRRRRRRNVsOR0RR:RR=FR50sEC#>R=R''42R;
RRRRRCRRDV#HRDPNHb8VGRR=b_F#xFCsRRFsPHND8GVbRM=RCxo_CRsF0MEC
RRRRRRRR-RR-CRs0MksRN#lD#DC0CR8MlFsNMDRkClLsR
RRRRRRRRR#MHoRRRRRR:=';j'
RRRRRRRRCRRGMbFRRRR:5=RFC0Es=#R>jR''
2;RRRRRRRRRsRVNRO0R:RR=FR50sEC#>R=R''j2R;
RRRRRRRRRNVsOj052=R:R''4;R
RRRRRRDRC#RHVPHND8GVbRb=RFM#_FNslDER0CRM
RRRRRRRRRRHVNRM85NVsOR02=4R''ER0CRMRR-RR-sRVNHO0FHMR#DRND4R""R3
RRRRRRRRRHRRVMRN8CR5GMbFRG5CbCFMMI0_HE80-84RF0IMF2R42RR='
4'RRRRRRRRRRRRRMRN8GRCbRFM5Rj2=jR''ER0CRM
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-GR bCFMMH0R#MRFCIRNNV$RsRFlHHMVM$H03R
RRRRRRRRRRRRRNC##sh0Rmq_W)hhQtR
RRRRRRRRRRRRRRCRsb0FsRmwpqta_ )h QuB_iHt'MN#0M_OCMCNl
RRRRRRRRRRRRRRRR"&Rwhu_ qXaw)a :CRhGV0q0RCsFsPCVIDF"R
RRRRRRRRRRRRRRCR#PHCs0I$RNHsMM
o;RRRRRRRRRRRRRCRs0MksR#bF_VHMV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRCFGbM=R:RbCGF+MRR
4;RRRRRRRRRRRRRsRVNRO0:5=RFC0Es=#R>jR''
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRDRC#RC
RRRRRRRRRVRRs0NORR:=VOsN0RR+4R;
RRRRRRRRR8CMR;HV
RRRRRRRR#CDHPVRN8DHVRbG=FRb#C_8MlFsN0DRE
CMRRRRRRRRRVRHR8NMRs5VN2O0R'=R40'RERCMRRRR-V-Rs0NOHRFMHN#RD"DR4
"3RRRRRRRRRRRR-s-RCs0kMlR#NCDD#b0RFH##LRDCMlFsNMDRkClLsR
RRRRRRRRRRGRCbRFMR:RR=FR50sEC#>R=R''j2R;
RRRRRRRRRCRRGMbF5Rj2:'=R4
';RRRRRRRRRRRRVOsN0RRRRR:=5EF0CRs#='>Rj;'2
RRRRRRRRCRRD
#CRRRRRRRRRRRRVOsN0=R:RNVsO+0RR
4;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVPHND8GVbRM=RCMo_FNslDER0CRM
RRRRRRRRRRHVF5sRVOsN0=2RR''jRC0EMRRRR-RR-sRVNHO0FHMR#DRNDjR""R3
RRRRRRRRRHRRVsRFRG5CbRFM5bCGFMMC0H_I8-0E4FR8IFM0R242R'=RjN'RMR8
RRRRRRRRRRRRRbCGF5MRj=2RR''4RC0EMRRRR-RR-lR1NCDD#C0RGMbFC
M0RRRRRRRRRRRRR-R-R0sCkRsM0RECDoNsCR#0MNCo0CHPRM8CFNslDkRMlsLC
RRRRRRRRRRRRCRRGMbFRR:=5EF0CRs#='>Rj;'2
RRRRRRRRRRRRVRRs0NORR:=5EF0CRs#='>R4;'2
RRRRRRRRRRRR#CDCR
RRRRRRRRRRRRRCFGbM=R:RbCGF-MRR
4;RRRRRRRRRRRRRsRVNRO0:5=RFC0Es=#R>4R''
2;RRRRRRRRRRRRCRM8H
V;RRRRRRRRRDRC#RC
RRRRRRRRRVRRs0NORR:=VOsN0RR-4R;
RRRRRRRRR8CMR;HV
RRRRRRRR#CDHPVRN8DHVRbG=CRMoC_8MlFsN0DRE
CMRRRRRRRRRVRHRRFs5NVsOV05s0NO'oEHEFR8IFM0R242R'=RjR'
RRRRRRRRRNRRMV8Rs0NOR25jR'=R40'RERCMR-RR-lR1NCDD#b0RFH##LRDCVOsN0MHF
RRRRRRRRRRRR0sCkRsMxFCsV5bRVOsN0MHF_8IH0=ER>sRVNHO0FIM_HE80,R
RRRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=C>RGMbFC_M0I0H8E
2;RRRRRRRRRDRC#RC
RRRRRRRRRVRRs0NORR:=VOsN0RR-4R;
RRRRRRRRR8CMR;HV
RRRRRRRR8CMR;HV
RRRRCRRD
#CRRRRRRRR-7-RCCOsNR#C0RECMLklCRs
RRRRRHRRVNRPDVH8b=GRR#bF_VHMRC0EMR
RRRRRRRRR-s-RCs0kMFRl#b0RF0#HHRPCMLklCRs
RRRRRRRRRbCGFRMRR:RR=FR50sEC#>R=R''42R;
RRRRRRRRRbCGF5MRj:2R=jR''R;
RRRRRRRRRNVsOR0RR:RR=FR50sEC#>R=R''42R;
RRRRRCRRDV#HRDPNHb8VGRR=b_F#xFCs
RRRRRRRRFRRsDRONV##bGR52RR=M_CoxFCsRC0EMR
RRRRRRRRR-s-RCs0kMlR#NCDD#M0RC0oNHRPC8FCMsDlNRlMkL
CsRRRRRRRRRHR#oRMRR:RR=4R''R;
RRRRRRRRRbCGFRMRR=R:R05FE#CsRR=>'2j';R
RRRRRRRRRVOsN0RRRRR:=5EF0CRs#='>Rj;'2
RRRRRRRRVRRs0NO5Rj2:'=R4
';RRRRRRRRCHD#VNRPDVH8b=GRRoMC_sMFlRND0MEC
RRRRRRRRHRRVMRN8VR5s0NO2RR='R4'0MECRRRRRR--VOsN0MHFRRH#NRDD"34"
RRRRRRRRRRRRRHVNRM85bCGF5MRCFGbM0CM_8IH04E-RI8FMR0F4R22=4R''R
RRRRRRRRRRRRRNRM8CFGbMjR52RR='Rj'0MEC
RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-- FGbM0CMRRH#FRMCN$INRFVslMRHVHHM0
$3RRRRRRRRRRRRR#RN#0CsR_hmWhq)Q
htRRRRRRRRRRRRRRRRsFCbsw0Rpamq_ht  B)Q_tui'#HM0ONMCN_MlRC
RRRRRRRRRRRRR&RRRu"w_Xh aaqw R):h0CGqCV0sPRFCDsVF
I"RRRRRRRRRRRRRRRR#CCPs$H0RsINMoHM;R
RRRRRRRRRRRRRskC0sMMRCHo_MbVVRs5VNHO0FIM_HE80RR=>VOsN0MHF_8IH0
E,RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>GRCbCFMMI0_HE802R;
RRRRRRRRRCRRD
#CRRRRRRRRRRRRRGRCbRFM:C=RGMbFR4+R;RRRRRRR-w-Rs0NOHRFMFsPCVIDF
RRRRRRRRRRRRVRRs0NORR:=5EF0CRs#='>Rj;'2
RRRRRRRRRRRR8CMR;HV
RRRRRRRRCRRD
#CRRRRRRRRRRRRVOsN0=R:RNVsO+0RR
4;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVPHND8GVbRM=RC8o_CsMFlRND0MEC
RRRRRRRRHRRVMRN8VR5s0NO2RR='R4'0MECRRRRRR--VOsN0MHFRRH#NRDD"34"
RRRRRRRRRRRRR--skC0s#MRlDNDCR#0b#F#HCLDRsMFlRNDMLklCRs
RRRRRRRRRCRRGMbFRRRR:5=RFC0Es=#R>jR''
2;RRRRRRRRRRRRCFGbM25jRR:=';4'
RRRRRRRRRRRRNVsOR0RR=R:R05FE#CsRR=>'2j';R
RRRRRRRRRCCD#
RRRRRRRRRRRRNVsO:0R=sRVNRO0+;R4
RRRRRRRRCRRMH8RVR;
RRRRRCRRDV#HRDPNHb8VGRR=b_F#MlFsN0DRE
CMRRRRRRRRRVRHRRFs5NVsOR02=jR''ER0CRMRRRRR-V-Rs0NOHRFMHN#RD"DRj
"3RRRRRRRRRRRRHFVRsCR5GMbFRG5CbCFMMI0_HE80-84RF0IMF2R42RR='Rj'N
M8RRRRRRRRRRRRRGRCbRFM5Rj2=4R''ER0CRMRRRRR-1-RlDNDCR#0CFGbM0CM
RRRRRRRRRRRR-RR-CRs0MksRC0ERsDNo0C#R#bFHP0HCCR8MlFsNMDRkClLsR
RRRRRRRRRRRRRCFGbM=R:R05FE#CsRR=>'2j';R
RRRRRRRRRRRRRVOsN0=R:R05FE#CsRR=>'24';R
RRRRRRRRRRDRC#RC
RRRRRRRRRRRRRbCGF:MR=GRCbRFM-;R4
RRRRRRRRRRRRVRRs0NORR:=5EF0CRs#='>R4;'2
RRRRRRRRRRRR8CMR;HV
RRRRRRRRCRRD
#CRRRRRRRRRRRRVOsN0=R:RNVsO-0RR
4;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVPHND8GVbRb=RF8#_CsMFlRND0MEC
RRRRRRRRHRRVsRFRs5VN5O0VOsN0H'Eo8ERF0IMF2R42RR='
j'RRRRRRRRRRRRNRM8VOsN0jR52RR='R4'0MECRRRR-1-RlDNDCR#0b#F#HCLDRNVsOF0HMR
RRRRRRRRRRCRs0MksRsxCFRVb5NVsOF0HMH_I8R0E=V>Rs0NOH_FMI0H8ER,
RRRRRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>CFGbM0CM_8IH0;E2
RRRRRRRRCRRD
#CRRRRRRRRRRRRVOsN0=R:RNVsO-0RR
4;RRRRRRRRRMRC8VRH;R
RRRRRRMRC8VRH;R
RRRRRCRM8H
V;RRRRRCRs#0kDR45-RI8FMR0F-NVsOF0HMH_I820ER=R:R)zh p1me_ 7VNDF0s5VN2O0;R
RRRRRskC#D50RCFGbM0CM_8IH0-ER4FR8IFM0RRj2:z=Rh1) m pe7D_VF5N0CFGbM
2;RRRRRCRs#0kDRG5CbCFMMI0_HE802RRRRRRRRRRRR=R:Ro#HMR;
RRRRR0sCkRsMskC#D
0;RRRRCRM8H
V;RMRC8kRVMHO0FhMRCNG0Vs0C;R

RR--)kC0sRM#aCskRRHVX#RHRFkMss8CCI8RHR0EYR3
RMVkOF0HMMRzFCs8sRC85R
RR,RGR:$RR)zh p1me_ 7VNDF0R2RRRRRRRRRR-R-RFVDNM0HoFRbHRM0HkMb0R
RRCRs0MksRmAmph q
HRR#R
RRNRPsLHNDDCRV$b0bRC,s0Vb$RbC:NRPD_H8V0b#N;0C
LRRCMoH
RRRRbDV0C$bRR:=O#DN#RVb5;G2
RRRRbsV0C$bRR:=O#DN#RVb5;$2
RRRRRHV5bDV0C$bRM=RNFMRsVRDbb0$CRR=JCkH0N_MMsRF
RRRRRRRRbsV0C$bRM=RNFMRsVRsbb0$CRR=JCkH0N_MMsRF
RRRRRRRRbDV0C$bRH=R#FGRsVRsbb0$CRR=H2#GRC0EMR
RRRRRskC0s0MRs;kC
RRRR#CDCR
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RCRM8VOkM0MHFRFzMss8CC
8;
VRRk0MOHRFMwHHM05CR
RRRR:GRR)zh p1me_ 7VNDF0R2
RsRRCs0kMmRAmqp hR
RHR#
RPRRNNsHLRDCV#b_0CN0RP:RN8DH_#Vb0CN0;-RR-bRVRN#00RC
RoLCHRM
RVRRb0_#NR0C:B=RD#N#V5bRG
2;RRRRH5VRV#b_0CN0Rb=RFH#_MRV2F5sRV#b_0CN0RM=RCHo_MRV20MEC
RRRRsRRCs0kMsR0k
C;RRRRCCD#
RRRRsRRCs0kMNRVD;#C
RRRR8CMR;HV
CRRMV8Rk0MOHRFMwHHM0
C;
VRRk0MOHRFMQN#MM
R5RRRRGRR:z h)1emp V7_D0FN2R
RRCRs0MksRmAmph q
HRR#R
RRNRPsLHNDVCRb0_#NR0C:NRPD_H8V0b#N;0CR-R-RRVb#00NCR
RLHCoMR
RRbRV_N#00:CR=DRBNV##bGR52R;
RHRRVVR5b0_#NR0C=NRMMF2RsVR5b0_#NR0C=kRJH_C0M2NMRC0EMR
RRRRRskC0s0MRs;kC
RRRR#CDCR
RRRRRskC0sVMRNCD#;R
RRMRC8VRH;R
RCRM8VOkM0MHFRMQ#N
M;
-RR-kRwMHO0F0MRFCRs0MksRMOF#M0N0
#3RkRVMHO0FxMRCVsFb
R5RRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;R-C-RGMbFC
M0RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RFVDNV0_s0NOH_FMI0H8ER2R-V-Rs0NOH
FMRRRRskC0szMRh1) m pe7D_VF
N0R#RH
RRRRMOF#M0N0CRs#0kDRz:Rh1) m pe7D_VFRN05bCGFMMC0H_I8R0E8MFI0-FRVOsN0MHF_8IH0RE2:R=
RRRRR05FE#CsRR=>'2j';RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-RR-CRxsRF
RoLCHRM
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRsxCF;Vb
R
RVOkM0MHFRMMNV5bR
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq:pR=DRVF_N0CFGbM0CM_8IH0RE;RR--CFGbM0CM
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=DRVF_N0VOsN0MHF_8IH0RE2RR--VOsN0MHF
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820ER
:=RRRRRFR50sEC#>R=R''j2R;RRRRRRRRRRRRRRRRR-x-RC
sFRCRLo
HMRRRRskC#D50RCFGbM0CM_8IH04E-RI8FMR0Fj:2R=FR50sEC#>R=R''42R;
R-RR-GR bCFMMN0RD"DR4R"
RsRRCD#k0-R54R2RRRRRRRRRRRRRRRRRRRRRR=R:R''4;-RR-1RvAVRFRNwsOF0HM4R""R
RR-R-R0hFCw:RsRFlWi3RERNM" Q  0R1NNM8s(8R6VcRFAsRHsMN$DRwFHN0MuoRF0HM"R
RR-R-RCaERV8HVCCsMROCLIC0CRCMNHR#oDMNHRMohRqhNRM8NkRJHRC0hRqhH0#RE
N0RRRR-0-REvCR1FARVER0CsRwNHO0FHMR#RRN"R4"HNMRRo1HMHNDMhoRqRh,NRM8HN#R
RRRRR--"Rj"HNMRRHJkCh0Rq
h3RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMNRMM;Vb
R
RVOkM0MHFRNJMMRVb5R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)Rqp:V=RD0FN_bCGFMMC0H_I8;0ER-R-RbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820ER-R-RNVsOF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802=R:
RRRR5RRFC0Es=#R>jR''R2;RRRRRRRRRRRRRRRRRR--xFCs
LRRCMoH
RRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>4R''
2;RRRR- -RGMbFCRM0NRDD"
4"RRRRskC#D50R-NVsOF0HMH_I820ERRRRRRRRR:RR=4R''R;R-p-R1FARVsRwNHO0F"MR4R"
R-RR-BR5F8kDRPENCCRLCNMRML$RH
02RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMMRJNbMV;R

RMVkOF0HMFRb#M_HVRVb5R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)Rqp:V=RD0FN_bCGFMMC0H_I8;0ER-R-RbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820ER-R-RNVsOF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802=R:
RRRR5RRFC0Es=#R>jR''R2;RRRRRRRRRRRRRRRRRR--xFCs
LRRCMoH
RRRR#sCkRD05bCGFMMC0H_I8-0E4FR8IFM0RRj2:5=RFC0Es=#R>4R''R2;RR-- FGbM0CMRDNDR""4
RRRR0sCkRsMskC#D
0;RMRC8kRVMHO0FbMRFH#_MbVV;R

RMVkOF0HMCRMoM_HVRVb5R
RRFROMN#0MC0RGMbFC_M0I0H8ERR:hzqa)Rqp:V=RD0FN_bCGFMMC0H_I8;0ER-R-RbCGFMMC0R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820ER-R-RNVsOF0HMR
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802=R:
RRRR5RRFC0Es=#R>jR''R2;RRRRRRRRRRRRRRRRRR--xFCs
LRRCMoH
RRRR#sCkRD05bCGFMMC0H_I8R0E8MFI0jFR2=R:R05FE#CsRR=>'24';-RR-FR0bHRL0N#RD"DR4R"
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRoMC_VHMV
b;
VRRk0MOHRFMM_CoxFCsV5bR
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq:pR=DRVF_N0CFGbM0CM_8IH0RE;RR--CFGbM0CM
RRRRMOF#M0N0sRVNHO0FIM_HE80Rh:Rq)azq:pR=DRVF_N0VOsN0MHF_8IH0RE2RR--VOsN0MHF
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820ER
:=RRRRRFR50sEC#>R=R''j2R;RRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRRR-x-RC
sFRCRLo
HMRRRRskC#D50RCFGbM0CM_8IH0RE2:'=R4
';RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMCRMoC_xsbFV;R

RR--#CHx_#sCRsPC#MHF#R
RVOkM0MHFRsxCFRVb5R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RsPNHDNLC#RHRDFM$#RkCFRVsHR#xoHM
RRRR0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sxMRCVsFb
R5RRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRNVsOF0HMH_I8R0E=->R#CHx_#sC'IDF2R;
R8CMRMVkOF0HMCRxsbFV;R

RMVkOF0HMNRMMRVb5R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RsPNHDNLC#RHRDFM$#RkCFRVsHR#xoHM
RRRR0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sMMRNbMVRR5
RRRRRbCGFMMC0H_I8R0E=#>RH_xCs'C#EEHo,R
RRRRRVOsN0MHF_8IH0=ER>#R-H_xCs'C#D2FI;R
RCRM8VOkM0MHFRMMNV
b;
VRRk0MOHRFMJMMNV5bR
RRRRx#HCC_s#RR:z h)1emp V7_D0FN2RRRRRRRRR--PHNsNCLDRRH#F$MDRCk#RsVFRx#HH
MoRRRRskC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kMMRJNbMVRR5
RRRRRbCGFMMC0H_I8R0E=#>RH_xCs'C#EEHo,R
RRRRRVOsN0MHF_8IH0=ER>#R-H_xCs'C#D2FI;R
RCRM8VOkM0MHFRNJMM;Vb
R
RVOkM0MHFR#bF_VHMV5bR
RRRRx#HCC_s#RR:z h)1emp V7_D0FN2RRRRRRRRR--PHNsNCLDRRH#F$MDRCk#RsVFRx#HH
MoRRRRskC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kMFRb#M_HVRVb5R
RRRRRCFGbM0CM_8IH0=ER>HR#xsC_CE#'H,oE
RRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F;I2
CRRMV8Rk0MOHRFMb_F#HVMVb
;
RkRVMHO0FMMRCHo_MbVVRR5
R#RRH_xCsRC#:hRz)m 1p7e _FVDNR02RRRRR-RR-NRPsLHNDHCR#MRFDk$R#VCRF#sRHMxHoR
RRCRs0MksR)zh p1me_ 7VNDF0#RH
LRRCMoH
RRRR0sCkRsMM_CoHVMVb
R5RRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRNVsOF0HMH_I8R0E=->R#CHx_#sC'IDF2R;
R8CMRMVkOF0HMCRMoM_HV;Vb
R
RVOkM0MHFRoMC_sxCFRVb5R
RRHR#xsC_C:#RR)zh p1me_ 7VNDF0R2RRRRRR-R-RsPNHDNLC#RHRDFM$#RkCFRVsHR#xoHM
RRRR0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sMMRCxo_CVsFb
R5RRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRNVsOF0HMH_I8R0E=->R#CHx_#sC'IDF2R;
R8CMRMVkOF0HMCRMoC_xsbFV;-

-NbsoRlN#0$MEHC##V_FV-
-RDs0_M#$0#ECHF#RV
V
R-R-RGaC0RHFVOkM0MHF#R
R-b-RkFsb#RC:I0sHCV#RD0FNR0HMFRRNDCHMRm5haO REoNMCL8RN0#C$2bC
0RR$RbCvgepb#DkRRH#5''z,XR''',RjR',',4'R''Z,WR''',RpR',',]'R''-,sRCs2Fs;R
R0C$bRNOEsM_H8CCG8$_L_pveg#RHRsNsN5$R1_a7ztpmQRB2FBVR]qq)B)a ;R
R0C$bRpvegM_H8CCG8$_L_NOEs#RHRsNsN5$RB)]qq Ba)F2RVaR17p_zmBtQ;R
R0C$bRpvegkbD#M_H8CCG8$_L_NOEs#RHRsNsN5$RB)]qq Ba)F2RVeRvpDgbk
#;
ORRF0M#NRM0huA1RRRRRRRRRB:R]qq)B)a RRRRRRRRRRRR:B=R]qq)B)a 'DPN5j4n2R;R-#-RbCNORNOEs0NOCRs
RMOF#M0N0eRvp0g_FE_ON:sRRNOEsM_H8CCG8$_L_pveg=R:RX"zjW4Zp"]-;R
RO#FM00NMRNOEsF_0_pvegRR:vgep_8HMC8GC__L$OsENR
:=RRRR5''zRR=>',z'R''XRR=>',X'R''jRR=>',j'R''4RR=>',4'R''ZRR=>',Z'
RRRRWR''>R=R''W,pR''>R=R''p,]R''>R=R''],-R''>R=R''-,0RFE#CsRR=>'2z';R
RO#FM00NMRNOEsF_0_pvegkbD#RR:vgepb#Dk_8HMC8GC__L$OsENR
:=RRRR5''zRR=>',z'R''XRR=>',X'R''jRR=>',j'R''4RR=>',4'R''ZRR=>',Z'
RRRRWR''>R=R''W,pR''>R=R''p,]R''>R=R''],-R''>R=R''-,0RFE#CsRR=>CFsss
2;
-RR-kRbs#bFC1:R	#HbRHIE0#CRbCNO
bRRsCFO8CksRH#	bE_IH#0CbCNORR5
RpRRRH:RM0FkRhpQ H2R#R
RRNRPsLHNDsCRCmN8	RR:Apmm ;qh
RRRRsPNHDNLCRRORRRRRB:R]qq)B)a ;R
RLHCoMR
RRERIHRDCp=R/RDMkDMRN83RpN'DDDoCM0/ER=RRjDbFF
RRRRHRRVpR53DND5R42=RR''sRFRNp3D4D52RR=huA1RRFspD3ND254R]=Ra02RE
CMRRRRRRRRs8CNR,5DRRO,s8CNm;	2
RRRRCRRD
#CRRRRRRRRC0GH;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RCRM8bOsFCs8kC	R#HIb_ECH0#ObNC
;
R-R-RsbkbCF#:ERBC#O	RC0ERMbkON0k0MHFRRHMNHRDMRC
RFbsOkC8sOCRE	CO_MbkON0k0MHFRR5
RNRRsRoRRH:RM1RRah)QtR;
RORRFMDFRF:RkA0Rm mpqRh;RRRRRRRRRRRRR-RR-ERaCRsCIRN#NFRODRFMH0MREDCRH
MCRRRR8RF0RRR:FRk0Apmm ;qhRRRRRRRRRRRRRRRR-a-RECCsR#INR8NRFH0RMER0CHRDMRC
RoRRFRF8RF:RkA0Rm mpqRh;RRRRRRRRRRRRR-RR-sRakHCRVMRCFEkoRNOEs0NOCRs#VMFk8R
RRERONRs#:MRHRaQh )t 2#RH
RRRRR-- lGNb#DC3pRRCDoNRbHMkR0#NRsC"jjjjjjj"",Rjjjj3jjj"",Rjj:jjj:jjR"
RNRRD#HNRsGNoRRRRRRRRRRRR1:Rah)Qt4R5RR0FN'soDoCM0RE2HN#RsRo;RR--lCN	RRH08MFI0sFRNCMo
RRRRsPNHDNLCORHFMDF,8RHF:0RRmAmph q;RRRRR--HCM0sDMN
RRRRsPNHDNLCRR[:hRQa  t)=R:RRj;RRRRRRRRRR--OsEN0#CsRNsC8R
RLHCoMR
RRFRoFR8RRR:=V#NDCR;
RHRROFFDM=R:RDVN#
C;RRRRH08FR:RR=NRVD;#C
RRRRsVFRHHRMRR40NFRsDo'C0MoEFRDFRb
RRRRRRHVGoNs5RH2=RR''sRFRsGNo25HRh=RAR1uFGsRN5soH=2RRR]aF[sRRO=RE#NsRC0EMR
RRRRRRGRCH
0;RRRRRDRC#RHVGoNs5RH2=:R''ER0CRM
RRRRRHRROFFDM=R:Rk0sCR;
RRRRR#CDHGVRN5soH=2RR''3RC0EMR
RRRRRR8RHF:0R=sR0k
C;RRRRRDRC#RHVGoNsR25HRR/='R_'0MEC
RRRRRRRR:[R=RR[+;R4
RRRRCRRMH8RVR;
RCRRMD8RF;Fb
RRRRRHV[RR=OsEN#ER0CRM
RRRRRFoF8=R:Rk0sCR;RRRRRRRRRRRRRRRRRR-RR-ERaCRsCNRsCCkMFoOERENNsO#0CRR0Fs8CN
RRRR8CMR;HV
RRRRDOFF:MR=ORHFMDF;R
RRVRHRFH80MRN8ORHFMDFRC0EMR
RRRRR8RF0:V=RNCD#;R
RRDRC#RC
RRRRR08FRR:=H08F;R
RRMRC8VRH;R
RCRM8bOsFCs8kCEROC_O	bOkM00kNH;FM
R
R-b-RkFsb#RC:1sCNO#ECRDNRHRMCVRFsN:R""MRN8CRsbODNCH#R0HRI0NERR""33R
RbOsFCs8kCHRVGF_ODRFM5R
RRsRNoRRR:MRHFRk01Qa)h
t;RRRROsEN#RR:HHMRMo0CCRs2HR#
RNRRD#HNRsGNoRRRRRRRRRRRR1:Rah)Qt4R5RR0FN'soDoCM0RE2HN#RsRo;RR--lCN	RRH08MFI0sFRNCMo
RRRRsPNHDNLCRR[:hRQa  t)=R:RRj;RRRRRRRRRR--OsEN0#CsRNsC8R
RLHCoMR
RRFRVsRRHH4MRRR0FN'soDoCM0DERF
FbRRRRRVRHRsGNo25HR'=RRF'RsNRGsHo52RR=huA1RRFsGoNs5RH2=aR]RRFs[RR>OsEN#ER0CRM
RRRRRCRRG;H0
RRRRCRRDV#HRsGNo25HR'=R:0'RE
CMRRRRRRRRGoNsR25HRR:=';3'
RRRRCRRDV#HRsGNoHR52=R/R''_RC0EMR
RRRRRRRR[:[=RR4+R;R
RRRRRCRM8H
V;RRRRCRM8DbFF;R
RCRM8bOsFCs8kCHRVGF_OD;FM
R
RbOsFCs8kC)RWQRa 5R
RRRRpRRRRRRRR:MRHFRk0p Qh;RRRRRRRRRRRR-RR-MRHbRk0DCHM
RRRRpeqzR RR:RRRRHMRzRRh1) m pe7D_VF;N0R-R-RFVDNM0HoFRbHRM0HkMb0R
RRzRK1waQQR 7:MRHRRRR1 Q7R=R:RosHE
0;RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RH
RRRRsPNHDNLCRR#RRRR:aR1)tQh504RFNRPD'kCEEHoRP-RNCDk'IDFR2+d;R
RRNRPsLHND#CRHGM8RQ:Rhta  
);RCRLoRHMRR--VOkM0MHFRHIs0RC
R#RR5R42RR:=vgep__0FOsEN571a_mzpt5QBezqp q5ep'z EEHo2;22
RRRR.#52:RR=:R''R;
R#RRHGM8RR:=dR;
RVRRFHsRRRHMezqp H'Eo4E-RI8FMR0FjFRDFRb
RRRRR##5HGM82=R:RpvegF_0_NOEsa517p_zmBtQ5peqzH 52;22
RRRR#RRHGM8RRRR:#=RHGM8R4+R;R
RRMRC8FRDF
b;RRRR#H5#M28GRR:=';:'
RRRRM#H8RGRR=R:RM#H8+GRR
4;RRRRVRFsHMRHRR-48MFI0eFRq pz'IDFRFDFbR
RRRRR#H5#M28GRR:=vgep__0FOsEN571a_mzpt5QBezqp 25H2
2;RRRRRHR#MR8GR:RR=HR#MR8G+;R4
RRRR8CMRFDFbR;
RWRR) QaR,5pRR#,Kaz1Q wQ7w,RQ7 p2R;
R8CMRFbsOkC8sWCR) Qa;R

RFbsOkC8s)CR Rq75:pRRFHMkp0RQ;h Rpeqz: RR0FkR)zh p1me_ 7VNDF0H2R#R
RR-R-R#uF#DHLCNR80RN:Rjj:j:jjjjjjj
jjRRRR-R-RRRRRRRRRRRRRRjRRjjjjjjjjj
jjRRRRPHNsNCLDRRORRRRR:]RBqB)qa; )
RRRRsPNHDNLCPRlRRRRRz:Rh1) m pe7D_VFRN05peqzs 'NCMo2R;
RPRRNNsHLRDCs8CNm:	RRmAmph q;R
RRNRPsLHNDDCRNk#0RRR:Apmm Rqh:V=RNCD#;RRRRRRRR-R-R#DN0ERONOsN0RCsIRN#N"MR_R"
RPRRNNsHLRDCHRRRR:RRRaQh )t ;RRRRRRRR-RR-MRH8RCGPHNsNCLD
LRRCMoHR-R-Rq) 7R
RRqRepRz :5=Rezqp N'sMRoC='>Rz;'2RRRRR-R-RHHM0DHNHRxC0NFRR""z
RRRRH1	bE_IH#0CbCNOR25p;R
RR R)q57RDO,R,CRsN	8m2R;
RHRRVqRep'z DoCM0>ERR0jRE
CMRRRRRRRH:P=RNCDk'oEHER;
RRRRRNsC8FDFbRR:DbFF
RRRRRRRRRHVs8CNm=	RRDVN#0CRERCMRRRRRRRRRR--ADNHR0FkRRHV0sECCNRI#RRNLRN8s8CN
RRRRRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCR
RRRRRRRRRRRR&"q) 7D5VF2N0:
R"RRRRRRRRRRRR& R"sssFR8CMRRFVVCHDROCMF0kMC8sC3R"
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCk;sM
RRRRRRRR#CDHOVRR'=RRF'RsRRO=)RBRRFsORR=]0aRERCMRR--s8CNHRMo8CFM3R
RRRRRRRRRH5VRH=R/RDPNkDC'FRI20MEC
RRRRRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRRRRRRRRR&"q) 7D5VF2N0:
R"RRRRRRRRRRRRRRR&"sWNMoHM:NReDRkC0MskOCN08
3"RRRRRRRRRRRRRCR#PHCs0I$RNHsMM
o;RRRRRRRRRRRRskC0s
M;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVORR='R_'0MEC
RRRRRRRRHRRVRRH=NRPD'kCEEHoRC0EMRRRRRRRRR--AHCoMI#RHR0EN"MR_R"
RRRRRRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCR
RRRRRRRRRRRRR&)R" 5q7VNDF0R2:"R
RRRRRRRRRRRRR&1R"0MsHoCRLo#HMR0IHEMRNR_"""R""#CCPs$H0RsCsF
s;RRRRRRRRRRRRskC0s
M;RRRRRRRRRDRC#RHVD0N#kER0CRMRRRRRRRRRRRRR-"-R_R_"8CC0O80C
RRRRRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_N
lCRRRRRRRRRRRRRRR&"q) 7D5VF2N0:
R"RRRRRRRRRRRRRRR&"FaIR8kMCOs#F#sCR08CCCO08MRHRbHMk#0R0MsHo"R"_"_""R
RRRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRRRRskC0s
M;RRRRRRRRRDRC#RC
RRRRRRRRRDRRNk#0RR:=0Csk;R
RRRRRRRRRCRM8H
V;RRRRRRRRCHD#VRRO=:R''sRFR=ORR''3RC0EMRRR-#-RCsbNNs0F,oRHMCFs
RRRRRRRRHRRVFRM0HR5R-=R4sRFR=HRRDPNkEC'H-oE402RE
CMRRRRRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_MlRC
RRRRRRRRRRRRR"&R)7 q5FVDN:02R
R"RRRRRRRRRRRRRRR&"sWNMoHM:CR1bNNs0RFsbMFH0FR8CM#RFl0RNE0ORlMkLRCsVlFsNR0:'R"
RRRRRRRRRRRRRO&RR"&R'MRCOMFk0CCs80RNRODFNF0HMRR"&hRQa  t)l'HN5oCH&2RR""3
RRRRRRRRRRRR#RRCsPCHR0$IMNsH;Mo
RRRRRRRRCRRMH8RVR;
RRRRRRRRR#DN0:kR=NRVD;#C
RRRRRRRR#CDH5VROsEN__0Fvgepb#Dk5RO2=sRCs2FsRC0EMR
RRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_MlRC
RRRRRRRRR&RRR ")qV75D0FN2":R
RRRRRRRRRRRR"&R FsssB:RENNsOs0CRR'"&RRO&'R"RNsC8C,RGObC0RC81_a7ztpmQDBRHs0CN"D3
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRD
#CRRRRRRRRRPRlR25HRR:=OsEN__0Fvgep5;O2
RRRRRRRRHRRRR:=HRR-4R;
RRRRRRRRRRHVHRR<PkNDCF'DIER0CRM
RRRRRRRRReRRq pzRR:=l
P;RRRRRRRRRRRRskC0s
M;RRRRRRRRRMRC8VRH;R
RRRRRRRRRD0N#k=R:RDVN#
C;RRRRRRRRCRM8H
V;RRRRRRRR)7 qR,5DRRO,s8CNm;	2
RRRRCRRMD8RFRFbs8CNDbFF;R
RRMRC8VRH;R
RCRM8bOsFCs8kC R)q
7;
bRRsCFO8CksRq) 7pR5RH:RM0FkRhpQ e;Rq pzRF:Rkz0Rh1) m pe7D_VF;N0Rmtm7RR:FRk0Apmm 2qhR
H#RRRR-u-RFH##LRDC8NN0:jRR:jjjjj:jjjjjjR
RR-R-RRRRRRRRRRRRRRRRRjjjjjjjjjjjjR
RRNRPsLHNDOCRRRRRRRR:B)]qq Ba)R;
RPRRNNsHLRDClRPRR:RRR)zh p1me_ 7VNDF0eR5q pz'MsNo;C2
RRRRsPNHDNLCNRD#R0kRA:Rm mpq:hR=NRVD;#CRRRRRRRRRR--D0N#RNOEs0NOCIsRNN#RM_R""R
RRNRPsLHNDHCRRRRRRRR:Q hat; )RRRRRRRRR-R-R8HMCPGRNNsHL
DCRRRRPHNsNCLDRNsC8Rm	:mRAmqp hR;
RoLCHRMR-)-R 
q7RRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;RRRRR-H-RMHH0NxDHCFR0R"NRzR"
R1RR	_HbI0EHCN#bO5CRp
2;RRRR)7 qR,5DRRO,s8CNm;	2
RRRRRHVezqp C'DMEo0Rj>RRC0EMR
RRRRRH=R:RDPNkEC'H;oE
RRRRoRRFRF8:V=RNCD#;R
RRRRRs8CNDbFFRD:RF
FbRRRRRRRRHsVRCmN8	RR=V#NDCER0CRMRRRRRRRRR-A-RNRHDFRk0H0VRECCsR#INRLNRNs8RC
N8RRRRRRRRRCRs0Mks;R
RRRRRRDRC#RHVORR='RR'FOsRRB=R)sRFR=ORRR]a0MECR-R-RNsC8oHMRM8FCR
RRRRRRRRRskC0s
M;RRRRRRRRCHD#VRRO=_R''ER0CRM
RRRRRRRRRRHVHRR=jER0CRMRRRRRRRRRRRRRR-RR-CRAo#HMR0IHEMRNR""_
RRRRRRRRRRRR0sCk;sM
RRRRRRRRCRRDV#HR#DN00kRERCMRRRRRRRRRRRRRR--""__R08CCCO08R
RRRRRRRRRRCRs0Mks;R
RRRRRRRRRCCD#
RRRRRRRRRRRR#DN0:kR=sR0k
C;RRRRRRRRRMRC8VRH;R
RRRRRRDRC#RHVORR='R:'FOsRR'=R30'RERCMR-R-Rb#CN0sNFRs,HFoMsRC
RRRRRRRRRR--o8FFRR:=5=HRRR-4FHsRRP=RNCDk'oEHE2-4;R
RRRRRRRRRD0N#k=R:RDVN#
C;RRRRRRRRCHD#VOR5E_Ns0vF_ebpgD5k#O=2RRsCsFRs20MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRD
#CRRRRRRRRRPRlR25HRR:=OsEN__0Fvgep5;O2
RRRRRRRRHRRRR:=HRR-4R;
RRRRRRRRRRHVHRR<PkNDCF'DIER0CRM
RRRRRRRRRoRRFRF8RR:=0Csk;R
RRRRRRRRRRqRepRz :l=RPR;
RRRRRRRRRsRRCs0kMR;
RRRRRRRRR8CMR;HV
RRRRRRRRDRRNk#0RR:=V#NDCR;
RRRRRCRRMH8RVR;
RRRRR)RR Rq75RD,Os,RCmN8	
2;RRRRRMRC8FRDFsbRCDN8F;Fb
RRRR#CDCR
RRRRRo8FFRR:=0Csk;RRRRRRRRRRRRRRRRRRRR-R-RNsC8MRH0NFRRDMkDsRNs
N$RRRRCRM8H
V;RMRC8sRbF8OCkRsC)7 q;R

RFbsOkC8smCRWa)Q 
R5RRRRpRRRRRRRRRR:HkMF0QRphR ;RRRRRRRRRRRRRR--NCOO#0#R$RbC5HbFMs0C2R
RRqRepRz RRRR:MRHRRRRz h)1emp V7_D0FN;-RR-NRPDRkC0IFRsCH0
RRRR1KzaQQw :7RRRHMR1RRQR7 RR:=sEHo0R;RR-R-RHIEO#ERHR8C0[FRkH#0V0$RC
G0RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RHRRRRRR--I0H8EVRFRCVHDR8
RoLCHRM
RWRR) QaRR5pRRRRRRRR=p>R,R
RRRRRRRRRRpeqzR RR=RR>FR0_0F#soHM5peqz, 2
RRRRRRRRRRRKaz1Q wQ7>R=R1KzaQQw 
7,RRRRRRRRRwRRQ7 pRRRRRR=>wpQ 7
2;RMRC8sRbF8OCkRsCmQW)a
 ;
bRRsCFO8CksR m)q57RpRR:HkMF0QRphR ;ezqp RR:FRk0z h)1emp V7_D0FN2#RH
RRRRMOF#M0N0CRMRRRRRRRRRQ:Rhta  :)R=5R5PkNDCC'DMEo0+/.2d*2RRRd;R-R-R8bN
RRRRsPNHDNLCDR#PRRRRRRRR1:Rap7_mBtQ_Be aRm)5-MC4FR8IFM0R;j2RRRRR-R-RP#D
RRRRsPNHDNLCDR#PRkRRRRRRk:RVCHG8eR5q pz'MsNo;C2R-R-R#zMHCoM8HRVGRC8bMFH0R
RRNRPsLHNDOCRRRRRRRRRRRR:B)]qq Ba)R;
RPRRNNsHLRDCFR	RRRRRR:RRRmAmph q;R
RRNRPsLHNDMCR$DLLCRRRRRR:1_a7pQmtB _eB)amRR5.8MFI0jFR2R;RRRRRR-RR-RRdL#H0
RRRRsPNHDNLCFROD,FMR08FRA:Rm mpq
h;RCRLo
HMRRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;RRRRR-H-RMHH0NxDHCFR0R"NRzR"
R1RR	_HbI0EHCN#bO5CRp
2;RRRRHeVRq pz'MDCoR0E>RRj0MEC
RRRRORRE	CO_MbkON0k0MHFRs5NoRRR=p>R3DND,R
RRRRRRRRRRRRRRRRRRRRRRORRFMDFRR=>OFFDMR,
RRRRRRRRRRRRRRRRRRRRRRRR8RF0R>R=R08F,R
RRRRRRRRRRRRRRRRRRRRRRoRRFRF8RR=>F
	,RRRRRRRRRRRRRRRRRRRRRRRRRNOEs=#R>CRM/;d2
RRRRHRRVFRM0	RFRC0EMR
RRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNlR"&Rmq) 7":R
RRRRRRRR&RRRE"#FRs0#H0sMCoRMkOFM80C:RR"&3RpN
DDRRRRRRRRRRR&"CRMCR8#0EFRNRPC"RR&HCM0o'CsHolNCMR5C2/d
RRRRRRRR&RRRP"RN8DHR0FONODRENNsOs0C#
3"RRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRCRs0Mks;R
RRRRRCHD#VFR80ER0CRM
RRRRRmRR)7 qR,5pRP#DkF,R	R2;RRRRRRRRR-RR-CRsNH8R0HRD	NCRRQzwXR 7MLklCRs
RRRRRHRRVFRM0	RFRC0EMR
RRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_Ml&CRR)"m :q7RR"
RRRRRRRRR&RRRs"CsRFsCFMOkCM08CRsNM8HoaR1)tQhR&"RRNp3DRD
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCk;sM
RRRRRRRR#CDCR
RRRRRRRRRezqp =R:R)zh p1me_ 7VNDF0#R5D2Pk;R
RRRRRRMRC8VRH;R
RRRRRCHD#VFRODRFM0MEC
RRRRRRRR m)q57RpM,R$DLLCF,R	R2;RRRRRRRRRR--s8CNRC0ERo#HMHRL0R
RRRRRRVRHR0MFRRF	0MEC
RRRRRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCRR&" m)qR7:"R
RRRRRRRRRRRR&"8 MRRFV#H0sMCoRMkOFMs0CC
8"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0Mks;R
RRRRRRDRC#RHVML$LD5CR.FR8IFM0RR42/"=RjRj"0MEC
RRRRRRRRsRRCsbF0DRVF_N0oCCMs_HOb'	oH0M#NCMO_lMNCRR&" m)qR7:"R
RRRRRRRRRRRR&"DQDCDoNRo#HMHRL0aR1)tQhROCMF0kMC"8R
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RVR;
RRRRRsRRCRN85RD,OF,R	R2;RRRRRRRRRRRRR-RR-CRsN08REOCRFMDF
RRRRRRRRGVH_DOFF5MRpD3NDM,RC2/d;RRRRRRRR-R-RbsCDCNO#ER0CFRODRFMIEH0R"NR3
"3RRRRRRRRmq) 7pR5,DR#P5kR#kDP'oEHER-48MFI0#FRD'PkD2FI,	RF2R;R-s-RCRN8HD0RHR	CNwRzQ7X RlMkL
CsRRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_NRlC&mR")7 q:
R"RRRRRRRRRRRR&CR"sssFROCMF0kMCs8RCHN8M1oRah)QtRR"&3RpN
DDRRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0Mks;R
RRRRRRDRC#RC
RRRRRRRRRP#Dk#R5D'PkEEHo2=R:RLM$LRDC5;j2
RRRRRRRReRRq pzRR:=z h)1emp V7_D0FNRD5#P;k2
RRRRRRRR8CMR;HV
RRRRCRRD
#CRRRRRRRRmq) 7pR5,DR#PF,R	
2;RRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_NRlC&mR")7 q:
R"RRRRRRRRRRRR& R"sssFROCMF0kMC88RkMsHoCRsN
8"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0Mks;R
RRRRRRMRC8VRH;R
RRRRRRVRHRs5FRD5#PC5M-84RF0IMFqRep'z EEHo-peqzD 'F4I+2=2RR''42ER0CRM
RRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_NRlC&mR")7 q:
R"RRRRRRRRRRRR&eR"CFO0ssR0kNMO03C8"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s
M;RRRRRRRRCRM8H
V;RRRRRRRRezqp =R:R_0FVNDF0#R5DeP5q pz'oEHEq-ep'z DRFI8MFI0jFR2R,
RRRRRRRRRRRRRRRRRRRRRRRRRqRep'z EEHo,eR-q pz'IDF2R;
RRRRR8CMR;HV
RRRR8CMR;HV
CRRMb8RsCFO8CksR m)q
7;
bRRsCFO8CksR m)qp75RH:RM0FkRhpQ e;Rq pzRF:Rkz0Rh1) m pe7D_VF;N0Rmtm7RR:FRk0Apmm 2qhR
H#RRRRO#FM00NMRRMCRRRRRRRR:hRQa  t)=R:RP55NCDk'MDCo+0E.d2/2RR*dR;RRR--b
N8RRRRPHNsNCLDRP#DRRRRRRRR:aR17m_pt_QBea Bm5)RM4C-RI8FMR0FjR2;RRRRRR--#
DPRRRRPHNsNCLDRP#DkRRRRRRR:VRkH8GCRq5ep'z soNMCR2;RR--zHM#o8MCRGVHCb8RF0HM
RRRRsPNHDNLCRRORRRRRRRRRB:R]qq)B)a ;R
RRNRPsLHNDFCR	RRRRRRRRRR:Apmm ;qh
RRRRsPNHDNLC$RMLCLDRRRRR1:Rap7_mBtQ_Be aRm)58.RF0IMF2Rj;RRRRRRRR-R-RLdRH
0#RRRRPHNsNCLDRDOFFRM,8RF0:mRAmqp hR;
RoLCHRM
ReRRq pzRR:=5peqzs 'NCMoRR=>'2z';RRRR-RR-MRHHN0HDCHxRR0FNzR""R
RRmRtmR7R:V=RNCD#;R
RR	R1HIb_ECH0#ObNCpR52R;
RHRRVqRep'z DoCM0>ERR0jRE
CMRRRRREROC_O	bOkM00kNHRFM5oNsR=RR>3RpN,DD
RRRRRRRRRRRRRRRRRRRRRRRRFRODRFM=O>RFMDF,R
RRRRRRRRRRRRRRRRRRRRRR8RRFR0RRR=>8,F0
RRRRRRRRRRRRRRRRRRRRRRRRFRoFR8R=F>R	R,
RRRRRRRRRRRRRRRRRRRRRRRROsEN#>R=R/MCd
2;RRRRRVRHR0MFRRF	0MEC
RRRRRRRR0sCk;sM
RRRRCRRDV#HR08FRC0EMR
RRRRRR)Rm Rq75Rp,#kDP,	RF2R;RRRRRRRRRR-R-RNsC80RHR	DHCRRNzXwQ M7RkClLsR
RRRRRRVRHR0MFRRF	0MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRD
#CRRRRRRRRRqRepRz :z=Rh1) m pe7D_VFRN05P#Dk
2;RRRRRRRRCRM8H
V;RRRRRDRC#RHVOFFDMER0CRM
RRRRRmRR)7 qR,5pRLM$L,DCR2F	;RRRRRRRR-RR-CRsN08RE#CRHRoML
H0RRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRR0sCk;sM
RRRRRRRR#CDHMVR$DLLC.R5RI8FMR0F4/2R=jR"j0"RE
CMRRRRRRRRRCRs0Mks;R
RRRRRRMRC8VRH;R
RRRRRRCRsN58RDO,R,	RF2R;RRRRRRRRRRRRRR-R-RNsC8ER0CFROD
FMRRRRRRRRV_HGOFFDMpR53DND,CRM/;d2RRRRRRRRRR--sDCbN#OCRC0ERDOFFIMRHR0EN3R""R3
RRRRRmRR)7 qR,5pRP#Dk#R5D'PkEEHo-84RF0IMFDR#PDk'F,I2R2F	;-RR-CRsNH8R0HRD	NCRRQzwXR 7MLklCRs
RRRRRHRRVFRM0	RFRC0EMR
RRRRRRRRRskC0s
M;RRRRRRRRCCD#
RRRRRRRR#RRDRPk5P#DkH'EoRE2:M=R$DLLCjR52R;
RRRRRRRRRpeqz: R=hRz)m 1p7e _FVDN50R#kDP2R;
RRRRRCRRMH8RVR;
RRRRR#CDCR
RRRRRR)Rm Rq75Rp,#,DPR2F	;R
RRRRRRVRHR0MFRRF	0MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RVR;
RRRRRHRRVFR5s#R5DMP5CR-48MFI0eFRq pz'oEHEq-ep'z D+FI4R22=4R''02RE
CMRRRRRRRRRCRs0Mks;R
RRRRRRMRC8VRH;R
RRRRRRqRepRz :0=RFD_VFRN05P#D5peqzE 'H-oEezqp F'DIFR8IFM0R,j2
RRRRRRRRRRRRRRRRRRRRRRRRRRRezqp H'EoRE,-peqzD 'F;I2
RRRRCRRMH8RVR;
RRRRRmtm7=R:Rk0sCR;
RCRRMH8RVR;
R8CMRFbsOkC8smCR)7 q;R

RFbsOkC8s]CRWa)Q 
R5RRRRpRRRRRRRRRR:HkMF0QRphR ;RRRRRRRRRRRRRR--NCOO#0#R$RbC5HbFMs0C2R
RRqRepRz RRRR:MRHRRRRz h)1emp V7_D0FN;-RR-NRPDRkC0IFRsCH0
RRRR1KzaQQw :7RRRHMR1RRQR7 RR:=sEHo0R;RR-R-RHIEO#ERHR8C0[FRkH#0V0$RC
G0RRRRwpQ 7RRRRRR:HRMRRQRW7Ra]:j=R2#RHRRRRRR--I0H8EVRFRCVHDR8
RoLCHRM
RWRR) QaRR5pRRRRRRRR=p>R,R
RRRRRRRRRRpeqzR RR=RR>FR0_0E#soHM5peqz, 2
RRRRRRRRRRRKaz1Q wQ7>R=R1KzaQQw 
7,RRRRRRRRRwRRQ7 pRRRRRR=>wpQ 7
2;RMRC8sRbF8OCkRsC]QW)a
 ;
bRRsCFO8CksR ])q57RpRR:HkMF0QRphR ;ezqp RR:FRk0z h)1emp V7_D0FN2#RH
RRRRMOF#M0N0CRMRRRRRRRRRQ:Rhta  :)R=5R5PkNDCC'DMEo0+/d2c*2RRRc;R-R-R8bN
RRRRsPNHDNLCDR#PRRRRRRRR1:Rap7_mBtQ_Be aRm)5-MC4FR8IFM0R;j2RRRRR-R-RP#D
RRRRsPNHDNLCDR#PRkRRRRRRk:RVCHG8eR5q pz'MsNo;C2R-R-R#zMHCoM8HRVGRC8bMFH0R
RRNRPsLHNDOCRRRRRRRRRRRR:B)]qq Ba)R;
RPRRNNsHLRDCFR	RRRRRR:RRRmAmph q;R
RRNRPsLHNDMCR$DLLCRRRRRR:1_a7pQmtB _eB)amRR5d8MFI0jFR2R;RRRRRR-RR-RRcL#H0
RRRRsPNHDNLCFROD,FMR08FRA:Rm mpq
h;RCRLo
HMRRRRezqp =R:Rq5ep'z soNMC>R=R''z2R;RRRRR-H-RMHH0NxDHCFR0R"NRzR"
R1RR	_HbI0EHCN#bO5CRp
2;RRRRHeVRq pz'MDCoR0E>RRj0MEC
RRRRORRE	CO_MbkON0k0MHFRs5NoRRR=p>R3DND,R
RRRRRRRRRRRRRRRRRRRRRRORRFMDFRR=>OFFDMR,
RRRRRRRRRRRRRRRRRRRRRRRR8RF0R>R=R08F,R
RRRRRRRRRRRRRRRRRRRRRRoRRFRF8RR=>F
	,RRRRRRRRRRRRRRRRRRRRRRRRRNOEs=#R>CRM/;c2
RRRRHRRVFRM0	RFRC0EMR
RRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNlR"&R]q) 7":R
RRRRRRRR&RRRE"#FRs0#H0sMCoRMkOFM80C:RR"&3RpN
DDRRRRRRRRRRR&"CRMCR8#0EFRNRPC"RR&HCM0o'CsHolNCMR5C2/c
RRRRRRRR&RRRP"RN8DHRGECRNOEs0NOC3s#"R
RRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRskC0s
M;RRRRRDRC#RHV8RF00MEC
RRRRRRRR ])q57Rp#,RD,PkR2F	;RRRRRRRRRRRRR--s8CNRRH0DCH	RzNRw QX7kRMlsLC
RRRRRRRRRHVMRF0F0	RE
CMRRRRRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNlR"&R]q) 7":R
RRRRRRRRRRRR"&RCFsssMRCOMFk0RC8s8CNHRMo1Qa)h"tRRp&R3DND
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRD
#CRRRRRRRRRqRepRz :z=Rh1) m pe7D_VFRN05P#Dk
2;RRRRRRRRCRM8H
V;RRRRRDRC#RHVOFFDMER0CRM
RRRRR]RR)7 qR,5pRLM$L,DCR2F	;RRRRRRRR-RR-CRsN08RE#CRHRoML
H0RRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRRbsCFRs0VNDF0C_oMHCsO	_boM'H#M0NOMC_NRlC&]R")7 q:
R"RRRRRRRRRRRR& R"MF8RV0R#soHMROCMF0kMC8sC"R
RRRRRRRRRRCR#PHCs0C$RsssF;R
RRRRRRRRRskC0s
M;RRRRRRRRCHD#V$RMLCLDRR5d8MFI04FR2=R/Rj"jj0"RE
CMRRRRRRRRRCRsb0FsRFVDNo0_CsMCHbO_	Ho'MN#0M_OCMCNlR"&R]q) 7":R
RRRRRRRRRRRR"&RQCDDoRND#MHoR0LHR)1aQRhtCFMOkCM08
R"RRRRRRRRRRRR#CCPs$H0RsCsF
s;RRRRRRRRRCRs0Mks;R
RRRRRRMRC8VRH;R
RRRRRRCRsN58RDO,R,	RF2R;RRRRRRRRRRRRRR-R-RNsC8ER0CFROD
FMRRRRRRRRV_HGOFFDMpR53DND,CRM/;c2RRRRRRRRRR--sDCbN#OCRC0ERDOFFIMRHR0EN3R""R3
RRRRR]RR)7 qR,5pRP#Dk#R5D'PkEEHo-84RF0IMFDR#PDk'F,I2R2F	;-RR-CRsNH8R0HRD	NCRRQzwXR 7MLklCRs
RRRRRHRRVFRM0	RFRC0EMR
RRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_Ml&CRR)"] :q7RR"
RRRRRRRRR&RRRs"CsRFsCFMOkCM08CRsNM8HoaR1)tQhR&"RRNp3DRD
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCk;sM
RRRRRRRR#CDCR
RRRRRRRRR#kDPRD5#PEk'H2oERR:=ML$LD5CRj
2;RRRRRRRRRqRepRz :z=Rh1) m pe7D_VFRN05P#Dk
2;RRRRRRRRCRM8H
V;RRRRRDRC#RC
RRRRR]RR)7 qR,5pRP#D,	RF2R;
RRRRRHRRVFRM0	RFRC0EMR
RRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_Ml&CRR)"] :q7RR"
RRRRRRRRR&RRRs" sRFsCFMOkCM08kR8soHMRNsC8R"
RRRRRRRRR#RRCsPCHR0$CFsssR;
RRRRRRRRR0sCk;sM
RRRRRRRR8CMR;HV
RRRRRRRRRHV5RFs5P#D5-MC4FR8IFM0RpeqzE 'H-oEezqp F'DI2+42RR='24'RC0EMR
RRRRRRRRRsFCbsV0RD0FN_MoCCOsH_ob	'#HM0ONMCN_Ml&CRR)"] :q7RR"
RRRRRRRRR&RRRC"eOs0FRk0sM0ONC"83
RRRRRRRRRRRRP#CC0sH$sRCs;Fs
RRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RVR;
RRRRReRRq pzRR:=0VF_D0FNRD5#Pq5ep'z EEHo-peqzD 'F8IRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRpeqzE 'H,oERq-ep'z D2FI;R
RRRRRCRM8H
V;RRRRCRM8H
V;RMRC8sRbF8OCkRsC]q) 7
;
RsRbF8OCkRsC]q) 7pR5RH:RM0FkRhpQ e;Rq pzRF:Rkz0Rh1) m pe7D_VF;N0Rmtm7RR:FRk0Apmm 2qhR
H#RRRRO#FM00NMRRMCRRRRRRRR:hRQa  t)=R:RP55NCDk'MDCo+0Edc2/2RR*cR;RRR--b
N8RRRRPHNsNCLDRP#DRRRRRRRR:aR17m_pt_QBea Bm5)RM4C-RI8FMR0FjR2;RRRRRR--#
DPRRRRPHNsNCLDRP#DkRRRRRRR:VRkH8GCRq5ep'z soNMCR2;RR--zHM#o8MCRGVHCb8RF0HM
RRRRsPNHDNLCRRORRRRRRRRRB:R]qq)B)a ;R
RRNRPsLHNDFCR	RRRRRRRRRR:Apmm ;qh
RRRRsPNHDNLC$RMLCLDRRRRR1:Rap7_mBtQ_Be aRm)58dRF0IMF2Rj;RRRRRRRR-R-RLcRH
0#RRRRPHNsNCLDRDOFFRM,8RF0:mRAmqp hR;
RoLCHRM
ReRRq pzRR:=5peqzs 'NCMoRR=>'2z';RRRR-RR-MRHHN0HDCHxRR0FNzR""R
RRmRtmR7R:V=RNCD#;R
RR	R1HIb_ECH0#ObNCpR52R;
RHRRVqRep'z DoCM0>ERR0jRE
CMRRRRREROC_O	bOkM00kNHRFM5oNsR=RR>3RpN,DD
RRRRRRRRRRRRRRRRRRRRRRRRFRODRFM=O>RFMDF,R
RRRRRRRRRRRRRRRRRRRRRR8RRFR0RRR=>8,F0
RRRRRRRRRRRRRRRRRRRRRRRRFRoFR8R=F>R	R,
RRRRRRRRRRRRRRRRRRRRRRRROsEN#>R=R/MCc
2;RRRRRVRHR0MFRRF	0MEC
RRRRRRRR0sCk;sM
RRRRCRRDV#HR08FRC0EMR
RRRRRR)R] Rq75Rp,#kDP,	RF2R;RRRRRRRRRR-R-RNsC80RHR	DHCRRNzXwQ M7RkClLsR
RRRRRRVRHR0MFRRF	0MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRD
#CRRRRRRRRRqRepRz :z=Rh1) m pe7D_VFRN05P#Dk
2;RRRRRRRRCRM8H
V;RRRRRDRC#RHVOFFDMER0CRM
RRRRR]RR)7 qR,5pRLM$L,DCR2F	;RRRRRRRR-RR-CRsN08RE#CRHRoML
H0RRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRR0sCk;sM
RRRRRRRR#CDHMVR$DLLCdR5RI8FMR0F4/2R=jR"jRj"0MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RVR;
RRRRRsRRCRN85RD,OF,R	R2;RRRRRRRRRRRRR-RR-CRsN08REOCRFMDF
RRRRRRRRGVH_DOFF5MRpD3NDM,RC2/c;RRRRRRRR-R-RbsCDCNO#ER0CFRODRFMIEH0R"NR3
"3RRRRRRRR]q) 7pR5,DR#P5kR#kDP'oEHER-48MFI0#FRD'PkD2FI,	RF2R;R-s-RCRN8HD0RHR	CNwRzQ7X RlMkL
CsRRRRRRRRHMVRFF0R	ER0CRM
RRRRRRRRR0sCk;sM
RRRRRRRR#CDCR
RRRRRRRRR#kDPRD5#PEk'H2oERR:=ML$LD5CRj
2;RRRRRRRRRqRepRz :z=Rh1) m pe7D_VFRN05P#Dk
2;RRRRRRRRCRM8H
V;RRRRRDRC#RC
RRRRR]RR)7 qR,5pRP#D,	RF2R;
RRRRRHRRVFRM0	RFRC0EMR
RRRRRRRRRskC0s
M;RRRRRRRRCRM8H
V;RRRRRRRRH5VRF5sR#5DPM4C-RI8FMR0Fezqp H'EoeE-q pz'IDF+242R'=R4R'20MEC
RRRRRRRRsRRCs0kMR;
RRRRRCRRMH8RVR;
RRRRReRRq pzRR:=0VF_D0FNRD5#Pq5ep'z EEHo-peqzD 'F8IRF0IMF2Rj,R
RRRRRRRRRRRRRRRRRRRRRRRRRRpeqzE 'H,oERq-ep'z D2FI;R
RRRRRCRM8H
V;RRRRRmRtm:7R=sR0k
C;RRRRCRM8H
V;RMRC8sRbF8OCkRsC]q) 7
;
-s-R0#D_$EM0C##HR
FM-s-bNNolRM#$0#ECHF#_MR
RVOkM0MHFR_0F#H0sM5oRPkNDCRR:z h)1emp V7_D0FN2CRs0MksR)1aQRhtHR#
RPRRNNsHLRDC#RRRRRR:1Qa)h4t5RR0FPkNDCH'Eo-ERRDPNkDC'F+IRd
2;RRRRPHNsNCLDRM#H8:GRRaQh )t ;R
RLHCoM-RR-kRVMHO0FIMRsCH0
RRRR4#52:RR=eRvp0g_FE_ON1s5az7_pQmtBq5ep5z ezqp H'Eo2E22R;
R#RR5R.2RR:=';:'
RRRRM#H8:GR=;Rd
RRRRsVFRHHRMqRep'z EEHo-84RF0IMFRRjDbFF
RRRR#RR5M#H8RG2:v=Re_pg0OF_E5Ns1_a7ztpmQeB5q pz52H22R;
RRRRRM#H8RGRR=R:RM#H8+GRR
4;RRRRCRM8DbFF;R
RR5R##8HMG:2R=:R''R;
R#RRHGM8RRRR:#=RHGM8R4+R;R
RRFRVsRRHH-MR4FR8IFM0RpeqzD 'FDIRF
FbRRRRR5R##8HMG:2R=eRvp0g_FE_ON1s5az7_pQmtBq5ep5z H222;R
RRRRR#8HMGRRRRR:=#8HMGRR+4R;
RCRRMD8RF;Fb
RRRR0sCkRsM#R;
R8CMRMVkOF0HMFR0_s#0H;Mo
R
RVOkM0MHFR_0FEs#0HRMo5DPNk:CRR)zh p1me_ 7VNDF0s2RCs0kMaR1)tQhR
H#RRRRPHNsNCLDRP#DR1:Rap7_mBtQ_Be aRm)5DPNkDC'C0MoER-48MFI0jFR2R;
RoLCHRM
RVRRDbFFRV:RFHsRRRHM#'DPsoNMCFRDFRb
RRRRRP#D5RH2:0=RFj_X45ZRPkNDCR5H+NRPD'kCD2FI2R;
RCRRMD8RFRFbVFDFbR;
RsRRCs0kMFR0_0E#soHMRD5#P
2;RMRC8kRVMHO0F0MRF#_E0MsHo
;
RkRVMHO0F0MRF#_F0MsHoPR5NCDkRz:Rh1) m pe7D_VF2N0R0sCkRsM1Qa)hHtR#R
RRNRPsLHND#CRD:PRR71a_tpmQeB_ mBa)PR5NCDk'MDCo-0E4FR8IFM0R;j2
LRRCMoH
RRRRFVDF:bRRsVFRHHRMDR#PN'sMRoCDbFF
RRRR#RRDHP52=R:R_0FXZj4RN5PD5kCHRR+PkNDCF'DI;22
RRRR8CMRFDFbDRVF;Fb
RRRR0sCkRsM0FF_#H0sM5oR#2DP;R
RCRM8VOkM0MHFR_0FFs#0H;Mo
R
RVOkM0MHFRFVsl0_#soHMRR5
RLRR#H0sMRoRRRRRRRRRRRRRR:RRR)1aQ;htR-RR-HRLM$NsRs#0H
MoRRRRO#FM00NMRbCGFMMC0H_I8R0E:qRhaqz)p=R:RFVDNC0_GMbFC_M0I0H8ER;
RORRF0M#NRM0VOsN0MHF_8IH0:ERRahqzp)qRR:=VNDF0s_VNHO0FIM_HE802R
RRCRs0MksR)zh p1me_ 7VNDF0R
RHR#
RPRRNNsHLRDCskC#D:0RR)zh p1me_ 7VNDF0CR5GMbFC_M0I0H8EFR8IFM0Rs-VNHO0FIM_HE802R;
RPRRNNsHLRDCpRRRR:RRRhpQ R;
RPRRNNsHLRDCo8FFR:RRRmAmph q;R
RLHCoMR
RRRRp:M=RC1IRah)QtL'5#H0sM;o2
RRRRq) 7pR5,CRs#0kD,FRoF;82
RRRRN8CDODFNR0C5;p2
RRRR#N#CRs05FoF8R2
RRRRRbsCFRs0wqpma _thQ )Bi_utM'H#M0NOMC_N
lCRRRRRRR&"FVsl0_#soHM:NRA80R#soHMR&"RR0L#soHM
RRRR#RRCsPCHR0$CFsssR;
RsRRCs0kMCRs#0kD;R
RCRM8VOkM0MHFRFVsl0_#soHM;R

RMVkOF0HMsRVFFl_#H0sM5oR
RRRR0F#soHMRRRRRRRRRRRRRRRRR1:Rah)QtR;RRR--mNO0D0R#soHM
RRRRMOF#M0N0GRCbCFMMI0_HE80Rh:Rq)azq:pR=DRVF_N0CFGbM0CM_8IH0
E;RRRRO#FM00NMRNVsOF0HMH_I8R0E:qRhaqz)p=R:RFVDNV0_s0NOH_FMI0H8ER2
RsRRCs0kMhRz)m 1p7e _FVDNR0
R
H#RRRRPHNsNCLDR#sCkRD0:hRz)m 1p7e _FVDN50RCFGbM0CM_8IH08ERF0IMFVR-s0NOH_FMI0H8E
2;RRRRPHNsNCLDRRpRRRRR:QRph
 ;RRRRPHNsNCLDRFoF8RRR:mRAmqp hR;
RoLCHRM
RpRRRR:=MRCI1Qa)h5t'Fs#0H2Mo;R
RR)Rm Rq75Rp,skC#DR0,o8FF2R;
R8RRCDNDF0ONCpR52R;
RNRR#s#C0oR5F2F8
RRRRsRRCsbF0pRwm_qat  h)_QBu'itH0M#NCMO_lMNCR
RRRRR&VR"s_FlFs#0H:MoR8ANRs#0HRMo"RR&Fs#0H
MoRRRRRCR#PHCs0C$RsssF;R
RRCRs0MksR#sCk;D0
CRRMV8Rk0MOHRFMVlsF_0F#soHM;R

RMVkOF0HMsRVFEl_#H0sM5oR
RRRR0E#soHMRRRRRRRRRRRRRRRRR1:Rah)QtR;RRR--ERCG#H0sMRo
RORRF0M#NRM0CFGbM0CM_8IH0:ERRahqzp)qRR:=VNDF0G_CbCFMMI0_HE80;R
RRFROMN#0MV0Rs0NOH_FMI0H8ERR:hzqa)Rqp:V=RD0FN_NVsOF0HMH_I820E
RRRR0sCkRsMz h)1emp V7_D0FN
HRR#R
RRNRPsLHNDsCRCD#k0RR:z h)1emp V7_D0FNRG5CbCFMMI0_HE80RI8FMR0F-NVsOF0HMH_I820E;R
RRNRPsLHNDpCRRRRRRRR:p Qh;R
RRNRPsLHNDoCRFRF8RRR:Apmm ;qh
LRRCMoH
RRRR:pR=CRMIaR1)tQh'#5E0MsHo
2;RRRR]q) 7pR5,CRs#0kD,FRoF;82
RRRRN8CDODFNR0C5;p2
RRRR#N#CRs05FoF8R2
RRRRRbsCFRs0wqpma _thQ )Bi_utM'H#M0NOMC_N
lCRRRRRRR&"FVsl#_E0MsHoA:RN#8R0MsHoRR"&#RE0MsHoR
RRRRR#CCPs$H0RsCsF
s;RRRRskC0ssMRCD#k0R;
R8CMRMVkOF0HMsRVFEl_#H0sM
o;
VRRk0MOHRFMVlsF_s#0HRMo5R
RR#RL0MsHo:RRR)1aQ;htRRRRRRRRRRRRRRRRR-R-RMLHNRs$#H0sMRo
R#RRH_xCsRC#:hRz)m 1p7e _FVDNR02RRRRR-RR-#RkCV8RF#sRHMxHoMRFD
$RRRRRskC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kMsRVF#l_0MsHoLR5#H0sMRoRRRRRR>R=R0L#soHM,R
RRRRRRRRRRRRRRRRRRRRRRGRCbCFMMI0_HE80RR=>#CHx_#sC'oEHER,
RRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F;I2
CRRMV8Rk0MOHRFMVlsF_s#0H;Mo
R
RVOkM0MHFRFVsl#_F0MsHo
R5RRRRFs#0HRMoR1:Rah)QtR;RRRRRRRRRRRRRRRRR-m-ROD0NRs#0H
MoRRRR#CHx_#sCRz:Rh1) m pe7D_VF2N0RRRRRRRR-k-R#RC8VRFs#HHxMFoRMRD$
RRRR0sCkRsMz h)1emp V7_D0FNR
H#RCRLo
HMRRRRskC0sVMRs_FlFs#0HRMo50F#soHMRRRRRRRR=F>R#H0sM
o,RRRRRRRRRRRRRRRRRRRRRRRRRbCGFMMC0H_I8R0E=#>RH_xCs'C#EEHo,R
RRRRRRRRRRRRRRRRRRRRRRVRRs0NOH_FMI0H8E>R=RH-#xsC_CD#'F;I2
CRRMV8Rk0MOHRFMVlsF_0F#soHM;R

RMVkOF0HMsRVFEl_#H0sM5oR
RRRR0E#soHMRRR:1Qa)hRt;RRRRRRRRRRRRRRRRRR--ERCG#H0sMRo
R#RRH_xCsRC#:hRz)m 1p7e _FVDNR02RRRRR-RR-#RkCV8RF#sRHMxHoMRFD
$RRRRRskC0szMRh1) m pe7D_VFRN0HR#
RoLCHRM
RsRRCs0kMsRVFEl_#H0sM5oREs#0HRMoRRRRR=RR>#RE0MsHoR,
RRRRRRRRRRRRRRRRRRRRRRRRCFGbM0CM_8IH0=ER>HR#xsC_CE#'H,oE
RRRRRRRRRRRRRRRRRRRRRRRRsRVNHO0FIM_HE80RR=>-x#HCC_s#F'DI
2;RMRC8kRVMHO0FVMRs_FlEs#0H;Mo
M
C8NRbOo	NCFRL8V$RD0FN_MoCCOsH_ob	;